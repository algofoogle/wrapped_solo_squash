// This is the unpowered netlist.
module wrapped_solo_squash (active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input active;
 input wb_clk_i;
 input wb_rst_i;
 inout wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 inout [37:0] io_oeb;
 inout [37:0] io_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 inout [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire clknet_0_wb_clk_i;
 wire \adapter.blue ;
 wire \adapter.debug_design_reset ;
 wire \adapter.game.ballDirX ;
 wire \adapter.game.ballDirY ;
 wire \adapter.game.ballX[0] ;
 wire \adapter.game.ballX[1] ;
 wire \adapter.game.ballX[2] ;
 wire \adapter.game.ballX[3] ;
 wire \adapter.game.ballX[4] ;
 wire \adapter.game.ballX[5] ;
 wire \adapter.game.ballX[6] ;
 wire \adapter.game.ballX[7] ;
 wire \adapter.game.ballX[8] ;
 wire \adapter.game.ballY[0] ;
 wire \adapter.game.ballY[1] ;
 wire \adapter.game.ballY[2] ;
 wire \adapter.game.ballY[3] ;
 wire \adapter.game.ballY[4] ;
 wire \adapter.game.ballY[5] ;
 wire \adapter.game.ballY[6] ;
 wire \adapter.game.ballY[7] ;
 wire \adapter.game.green ;
 wire \adapter.game.h[0] ;
 wire \adapter.game.h[1] ;
 wire \adapter.game.h[2] ;
 wire \adapter.game.h[3] ;
 wire \adapter.game.h[4] ;
 wire \adapter.game.h[5] ;
 wire \adapter.game.h[6] ;
 wire \adapter.game.h[7] ;
 wire \adapter.game.h[8] ;
 wire \adapter.game.h[9] ;
 wire \adapter.game.hit ;
 wire \adapter.game.hsync ;
 wire \adapter.game.inBallX ;
 wire \adapter.game.inBallY ;
 wire \adapter.game.inPaddle ;
 wire \adapter.game.offset[0] ;
 wire \adapter.game.offset[1] ;
 wire \adapter.game.offset[2] ;
 wire \adapter.game.offset[3] ;
 wire \adapter.game.offset[4] ;
 wire \adapter.game.paddle[0] ;
 wire \adapter.game.paddle[1] ;
 wire \adapter.game.paddle[2] ;
 wire \adapter.game.paddle[3] ;
 wire \adapter.game.paddle[4] ;
 wire \adapter.game.paddle[5] ;
 wire \adapter.game.paddle[6] ;
 wire \adapter.game.paddle[7] ;
 wire \adapter.game.paddle[8] ;
 wire \adapter.game.red ;
 wire \adapter.game.speaker ;
 wire \adapter.game.v[0] ;
 wire \adapter.game.v[1] ;
 wire \adapter.game.v[2] ;
 wire \adapter.game.v[3] ;
 wire \adapter.game.v[4] ;
 wire \adapter.game.v[5] ;
 wire \adapter.game.v[6] ;
 wire \adapter.game.v[7] ;
 wire \adapter.game.v[8] ;
 wire \adapter.game.v[9] ;
 wire \adapter.game.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 sky130_fd_sc_hd__clkbuf_2 _0723_ (.A(net1),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_4 _0724_ (.A(_0057_),
    .X(_0058_));
 sky130_fd_sc_hd__inv_2 _0725_ (.A(_0058_),
    .Y(_0620_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(_0058_),
    .Y(_0621_));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(_0058_),
    .Y(_0622_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(_0058_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(_0058_),
    .Y(_0624_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(_0058_),
    .Y(_0625_));
 sky130_fd_sc_hd__buf_6 _0731_ (.A(_0057_),
    .X(_0059_));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(_0059_),
    .Y(_0626_));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(_0059_),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(_0059_),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(_0059_),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(_0059_),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(_0059_),
    .Y(_0523_));
 sky130_fd_sc_hd__buf_4 _0738_ (.A(_0057_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(_0060_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(_0060_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(_0060_),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(_0060_),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(_0060_),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(_0060_),
    .Y(_0529_));
 sky130_fd_sc_hd__buf_6 _0745_ (.A(_0057_),
    .X(_0061_));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(_0061_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(_0061_),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0061_),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(_0061_),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(_0061_),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(_0061_),
    .Y(_0535_));
 sky130_fd_sc_hd__clkbuf_4 _0752_ (.A(_0057_),
    .X(_0062_));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(_0062_),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0062_),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(_0062_),
    .Y(_0538_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(_0062_),
    .Y(_0539_));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(_0062_),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(_0062_),
    .Y(_0541_));
 sky130_fd_sc_hd__clkbuf_2 _0759_ (.A(net1),
    .X(_0063_));
 sky130_fd_sc_hd__buf_4 _0760_ (.A(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(_0064_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(_0064_),
    .Y(_0543_));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(_0064_),
    .Y(_0544_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(_0064_),
    .Y(_0545_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0064_),
    .Y(_0546_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(_0064_),
    .Y(_0547_));
 sky130_fd_sc_hd__buf_6 _0767_ (.A(_0063_),
    .X(_0065_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0065_),
    .Y(_0548_));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(_0065_),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0065_),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(_0065_),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(_0065_),
    .Y(_0553_));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(_0065_),
    .Y(_0554_));
 sky130_fd_sc_hd__buf_6 _0774_ (.A(_0063_),
    .X(_0066_));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(_0066_),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0066_),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(_0066_),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(_0066_),
    .Y(_0558_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(_0066_),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(_0066_),
    .Y(_0560_));
 sky130_fd_sc_hd__clkbuf_8 _0781_ (.A(_0063_),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(_0067_),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(_0067_),
    .Y(_0562_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(_0067_),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(_0067_),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(_0067_),
    .Y(_0565_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(_0067_),
    .Y(_0566_));
 sky130_fd_sc_hd__buf_4 _0788_ (.A(_0063_),
    .X(_0068_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(_0068_),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(_0068_),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(_0068_),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(_0068_),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(_0068_),
    .Y(_0572_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(_0068_),
    .Y(_0573_));
 sky130_fd_sc_hd__buf_4 _0795_ (.A(_0063_),
    .X(_0069_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(_0069_),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(_0069_),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(_0069_),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(_0069_),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(_0069_),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(_0069_),
    .Y(_0579_));
 sky130_fd_sc_hd__clkbuf_2 _0802_ (.A(net1),
    .X(_0070_));
 sky130_fd_sc_hd__buf_4 _0803_ (.A(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(_0071_),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(_0071_),
    .Y(_0581_));
 sky130_fd_sc_hd__inv_2 _0806_ (.A(_0071_),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(_0071_),
    .Y(_0583_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(_0071_),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(_0071_),
    .Y(_0585_));
 sky130_fd_sc_hd__buf_6 _0810_ (.A(_0070_),
    .X(_0072_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(_0072_),
    .Y(_0586_));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(_0072_),
    .Y(_0587_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(_0072_),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(_0072_),
    .Y(_0589_));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(_0072_),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(_0072_),
    .Y(_0592_));
 sky130_fd_sc_hd__clkbuf_8 _0817_ (.A(_0070_),
    .X(_0073_));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(_0073_),
    .Y(_0593_));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(_0073_),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(_0073_),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(_0073_),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(_0073_),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(_0073_),
    .Y(_0598_));
 sky130_fd_sc_hd__buf_4 _0824_ (.A(_0070_),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _0825_ (.A(_0074_),
    .Y(_0599_));
 sky130_fd_sc_hd__inv_2 _0826_ (.A(_0074_),
    .Y(_0600_));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(_0074_),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _0828_ (.A(_0074_),
    .Y(_0602_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(_0074_),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(_0074_),
    .Y(_0604_));
 sky130_fd_sc_hd__buf_4 _0831_ (.A(_0070_),
    .X(_0075_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(_0075_),
    .Y(_0605_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0075_),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _0834_ (.A(_0075_),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(_0075_),
    .Y(_0609_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(_0075_),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(_0075_),
    .Y(_0611_));
 sky130_fd_sc_hd__buf_6 _0838_ (.A(_0070_),
    .X(_0076_));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(_0076_),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_2 _0840_ (.A(_0076_),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0076_),
    .Y(_0614_));
 sky130_fd_sc_hd__inv_2 _0842_ (.A(_0076_),
    .Y(_0615_));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(_0076_),
    .Y(_0616_));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(_0076_),
    .Y(_0617_));
 sky130_fd_sc_hd__clkbuf_8 _0845_ (.A(net1),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _0846_ (.A(_0077_),
    .Y(_0618_));
 sky130_fd_sc_hd__inv_2 _0847_ (.A(_0077_),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _0848_ (.A(_0077_),
    .Y(_0608_));
 sky130_fd_sc_hd__inv_2 _0849_ (.A(_0077_),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _0850_ (.A(_0077_),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _0851_ (.A(_0077_),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _0852_ (.A(_0057_),
    .Y(_0519_));
 sky130_fd_sc_hd__and2b_1 _0853_ (.A_N(net7),
    .B(net5),
    .X(_0078_));
 sky130_fd_sc_hd__inv_2 _0854_ (.A(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0855_ (.A(_0079_),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _0856_ (.A(_0080_),
    .X(\adapter.debug_design_reset ));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(\adapter.game.h[7] ),
    .Y(_0081_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0858_ (.A(\adapter.game.h[5] ),
    .X(_0082_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0859_ (.A(\adapter.game.h[4] ),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_2 _0860_ (.A(\adapter.game.h[6] ),
    .X(_0084_));
 sky130_fd_sc_hd__nor3_1 _0861_ (.A(_0082_),
    .B(_0083_),
    .C(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__clkbuf_2 _0862_ (.A(\adapter.game.h[8] ),
    .X(_0086_));
 sky130_fd_sc_hd__a31o_1 _0863_ (.A1(_0082_),
    .A2(_0083_),
    .A3(_0084_),
    .B1(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_2 _0864_ (.A(\adapter.game.h[9] ),
    .X(_0088_));
 sky130_fd_sc_hd__or4b_1 _0865_ (.A(_0081_),
    .B(_0085_),
    .C(_0087_),
    .D_N(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_1 _0866_ (.A(_0089_),
    .X(\adapter.game.hsync ));
 sky130_fd_sc_hd__buf_2 _0867_ (.A(\adapter.game.v[9] ),
    .X(_0090_));
 sky130_fd_sc_hd__inv_2 _0868_ (.A(\adapter.game.v[3] ),
    .Y(_0091_));
 sky130_fd_sc_hd__clkbuf_2 _0869_ (.A(\adapter.game.v[2] ),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_2 _0870_ (.A(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_2 _0871_ (.A(\adapter.game.v[1] ),
    .X(_0094_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__or3_1 _0873_ (.A(_0091_),
    .B(_0093_),
    .C(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_2 _0874_ (.A(\adapter.game.v[4] ),
    .X(_0097_));
 sky130_fd_sc_hd__buf_2 _0875_ (.A(\adapter.game.v[8] ),
    .X(_0098_));
 sky130_fd_sc_hd__buf_2 _0876_ (.A(\adapter.game.v[7] ),
    .X(_0099_));
 sky130_fd_sc_hd__buf_2 _0877_ (.A(\adapter.game.v[5] ),
    .X(_0100_));
 sky130_fd_sc_hd__and4_1 _0878_ (.A(_0098_),
    .B(_0099_),
    .C(\adapter.game.v[6] ),
    .D(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__or4b_1 _0879_ (.A(_0090_),
    .B(_0096_),
    .C(_0097_),
    .D_N(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _0880_ (.A(_0102_),
    .X(\adapter.game.vsync ));
 sky130_fd_sc_hd__o21a_1 _0881_ (.A1(\adapter.game.h[7] ),
    .A2(_0086_),
    .B1(\adapter.game.h[9] ),
    .X(_0103_));
 sky130_fd_sc_hd__a31o_1 _0882_ (.A1(\adapter.game.h[5] ),
    .A2(_0084_),
    .A3(_0088_),
    .B1(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__a31o_1 _0883_ (.A1(\adapter.game.v[8] ),
    .A2(\adapter.game.v[7] ),
    .A3(\adapter.game.v[6] ),
    .B1(\adapter.game.v[9] ),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _0884_ (.A(\adapter.game.v[9] ),
    .B(\adapter.game.v[8] ),
    .X(_0106_));
 sky130_fd_sc_hd__or3_1 _0885_ (.A(\adapter.game.v[7] ),
    .B(\adapter.game.v[6] ),
    .C(\adapter.game.v[5] ),
    .X(_0107_));
 sky130_fd_sc_hd__nor2_1 _0886_ (.A(_0106_),
    .B(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__or3_1 _0887_ (.A(_0104_),
    .B(_0105_),
    .C(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__a21oi_1 _0888_ (.A1(\adapter.game.inBallY ),
    .A2(\adapter.game.inBallX ),
    .B1(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__nor3_1 _0889_ (.A(_0090_),
    .B(_0101_),
    .C(_0103_),
    .Y(_0111_));
 sky130_fd_sc_hd__and2b_1 _0890_ (.A_N(_0110_),
    .B(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0891_ (.A(_0112_),
    .X(\adapter.game.green ));
 sky130_fd_sc_hd__nor3_1 _0892_ (.A(\adapter.game.h[5] ),
    .B(\adapter.game.h[6] ),
    .C(\adapter.game.h[7] ),
    .Y(_0113_));
 sky130_fd_sc_hd__and4bb_1 _0893_ (.A_N(_0088_),
    .B_N(_0086_),
    .C(_0113_),
    .D(\adapter.game.inPaddle ),
    .X(_0114_));
 sky130_fd_sc_hd__or2_1 _0894_ (.A(\adapter.game.v[4] ),
    .B(\adapter.game.v[1] ),
    .X(_0115_));
 sky130_fd_sc_hd__nand2_1 _0895_ (.A(\adapter.game.v[3] ),
    .B(\adapter.game.v[2] ),
    .Y(_0116_));
 sky130_fd_sc_hd__o2bb2a_1 _0896_ (.A1_N(\adapter.game.v[4] ),
    .A2_N(_0094_),
    .B1(_0092_),
    .B2(\adapter.game.v[3] ),
    .X(_0117_));
 sky130_fd_sc_hd__a21oi_1 _0897_ (.A1(_0115_),
    .A2(_0116_),
    .B1(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__clkbuf_2 _0898_ (.A(\adapter.game.h[3] ),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_2 _0899_ (.A(\adapter.game.h[2] ),
    .X(_0120_));
 sky130_fd_sc_hd__and4_1 _0900_ (.A(\adapter.game.h[1] ),
    .B(_0119_),
    .C(_0120_),
    .D(\adapter.game.h[4] ),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_2 _0901_ (.A(\adapter.game.h[1] ),
    .X(_0122_));
 sky130_fd_sc_hd__nor4_1 _0902_ (.A(_0122_),
    .B(_0119_),
    .C(_0120_),
    .D(_0083_),
    .Y(_0123_));
 sky130_fd_sc_hd__o31a_1 _0903_ (.A1(_0118_),
    .A2(_0121_),
    .A3(_0123_),
    .B1(_0109_),
    .X(_0124_));
 sky130_fd_sc_hd__o21ai_2 _0904_ (.A1(_0114_),
    .A2(_0124_),
    .B1(_0111_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _0905_ (.A(_0125_),
    .Y(\adapter.game.red ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0906_ (.A(\adapter.game.ballY[6] ),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_2 _0907_ (.A(\adapter.game.ballY[5] ),
    .X(_0127_));
 sky130_fd_sc_hd__and2_1 _0908_ (.A(\adapter.game.ballY[3] ),
    .B(\adapter.game.ballY[4] ),
    .X(_0128_));
 sky130_fd_sc_hd__or2_1 _0909_ (.A(_0127_),
    .B(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0910_ (.A(\adapter.game.ballY[4] ),
    .X(_0130_));
 sky130_fd_sc_hd__nor4_1 _0911_ (.A(_0130_),
    .B(_0127_),
    .C(_0126_),
    .D(\adapter.game.ballY[7] ),
    .Y(_0131_));
 sky130_fd_sc_hd__clkbuf_2 _0912_ (.A(\adapter.game.ballX[6] ),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_2 _0913_ (.A(\adapter.game.ballX[7] ),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_2 _0914_ (.A(\adapter.game.ballX[3] ),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_2 _0915_ (.A(\adapter.game.ballX[4] ),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_2 _0916_ (.A(\adapter.game.ballX[5] ),
    .X(_0136_));
 sky130_fd_sc_hd__o21a_1 _0917_ (.A1(_0134_),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__o31a_1 _0918_ (.A1(_0132_),
    .A2(_0133_),
    .A3(_0137_),
    .B1(\adapter.game.ballX[8] ),
    .X(_0138_));
 sky130_fd_sc_hd__a311o_1 _0919_ (.A1(_0126_),
    .A2(\adapter.game.ballY[7] ),
    .A3(_0129_),
    .B1(_0131_),
    .C1(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_2 _0920_ (.A(\adapter.game.v[6] ),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _0921_ (.A1(_0100_),
    .A2(\adapter.game.hit ),
    .B1(_0139_),
    .B2(_0140_),
    .X(\adapter.game.speaker ));
 sky130_fd_sc_hd__inv_2 _0922_ (.A(\adapter.game.v[0] ),
    .Y(_0141_));
 sky130_fd_sc_hd__or2b_1 _0923_ (.A(\adapter.game.offset[2] ),
    .B_N(\adapter.game.v[1] ),
    .X(_0142_));
 sky130_fd_sc_hd__and2b_1 _0924_ (.A_N(\adapter.game.v[1] ),
    .B(\adapter.game.offset[2] ),
    .X(_0143_));
 sky130_fd_sc_hd__a31o_1 _0925_ (.A1(_0141_),
    .A2(\adapter.game.offset[1] ),
    .A3(_0142_),
    .B1(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0926_ (.A(\adapter.game.offset[2] ),
    .X(_0145_));
 sky130_fd_sc_hd__or2b_1 _0927_ (.A(\adapter.game.h[1] ),
    .B_N(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__or2b_1 _0928_ (.A(\adapter.game.h[0] ),
    .B_N(\adapter.game.offset[1] ),
    .X(_0147_));
 sky130_fd_sc_hd__and2b_1 _0929_ (.A_N(_0145_),
    .B(\adapter.game.h[1] ),
    .X(_0148_));
 sky130_fd_sc_hd__a21o_1 _0930_ (.A1(_0146_),
    .A2(_0147_),
    .B1(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__xnor2_1 _0931_ (.A(_0092_),
    .B(\adapter.game.h[2] ),
    .Y(_0150_));
 sky130_fd_sc_hd__xnor2_1 _0932_ (.A(_0149_),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__xnor2_1 _0933_ (.A(_0144_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(\adapter.game.offset[3] ),
    .Y(_0153_));
 sky130_fd_sc_hd__a221o_1 _0935_ (.A1(_0153_),
    .A2(\adapter.game.h[2] ),
    .B1(_0146_),
    .B2(_0147_),
    .C1(_0148_),
    .X(_0154_));
 sky130_fd_sc_hd__o21ai_1 _0936_ (.A1(_0153_),
    .A2(_0120_),
    .B1(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__and2b_1 _0937_ (.A_N(\adapter.game.offset[4] ),
    .B(\adapter.game.h[3] ),
    .X(_0156_));
 sky130_fd_sc_hd__and2b_1 _0938_ (.A_N(_0119_),
    .B(\adapter.game.offset[4] ),
    .X(_0157_));
 sky130_fd_sc_hd__nor2_1 _0939_ (.A(_0156_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__xnor2_1 _0940_ (.A(_0155_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_1 _0941_ (.A(_0092_),
    .B(_0153_),
    .Y(_0160_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(\adapter.game.v[2] ),
    .B(_0153_),
    .Y(_0161_));
 sky130_fd_sc_hd__a21oi_1 _0943_ (.A1(_0160_),
    .A2(_0144_),
    .B1(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__and2_1 _0944_ (.A(_0091_),
    .B(\adapter.game.offset[4] ),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_1 _0945_ (.A(_0091_),
    .B(\adapter.game.offset[4] ),
    .Y(_0164_));
 sky130_fd_sc_hd__nor2_1 _0946_ (.A(_0163_),
    .B(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__xnor2_1 _0947_ (.A(_0162_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__xnor2_1 _0948_ (.A(_0159_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__xnor2_1 _0949_ (.A(_0152_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__clkbuf_2 _0950_ (.A(\adapter.game.v[0] ),
    .X(_0169_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0951_ (.A(\adapter.game.h[0] ),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_1 _0952_ (.A(_0169_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__and2_1 _0953_ (.A(_0169_),
    .B(\adapter.game.h[0] ),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_1 _0954_ (.A(_0164_),
    .B(_0162_),
    .Y(_0173_));
 sky130_fd_sc_hd__or2_1 _0955_ (.A(_0163_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__or2b_1 _0956_ (.A(\adapter.game.offset[4] ),
    .B_N(_0119_),
    .X(_0175_));
 sky130_fd_sc_hd__a21oi_1 _0957_ (.A1(_0175_),
    .A2(_0155_),
    .B1(_0157_),
    .Y(_0176_));
 sky130_fd_sc_hd__xor2_1 _0958_ (.A(_0097_),
    .B(\adapter.game.h[4] ),
    .X(_0177_));
 sky130_fd_sc_hd__xnor2_1 _0959_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__xnor2_1 _0960_ (.A(_0174_),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__o31ai_1 _0961_ (.A1(_0168_),
    .A2(_0171_),
    .A3(_0172_),
    .B1(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__o211a_1 _0962_ (.A1(_0179_),
    .A2(_0168_),
    .B1(_0110_),
    .C1(_0125_),
    .X(_0181_));
 sky130_fd_sc_hd__and2b_1 _0963_ (.A_N(\adapter.game.offset[1] ),
    .B(_0172_),
    .X(_0182_));
 sky130_fd_sc_hd__a211o_1 _0964_ (.A1(\adapter.game.offset[1] ),
    .A2(_0171_),
    .B1(_0182_),
    .C1(_0179_),
    .X(_0183_));
 sky130_fd_sc_hd__and3_1 _0965_ (.A(_0180_),
    .B(_0181_),
    .C(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0966_ (.A(_0184_),
    .X(\adapter.blue ));
 sky130_fd_sc_hd__and2_1 _0967_ (.A(\adapter.game.h[9] ),
    .B(\adapter.game.h[8] ),
    .X(_0185_));
 sky130_fd_sc_hd__and4_1 _0968_ (.A(\adapter.game.h[1] ),
    .B(\adapter.game.h[0] ),
    .C(\adapter.game.h[3] ),
    .D(\adapter.game.h[2] ),
    .X(_0186_));
 sky130_fd_sc_hd__and4_1 _0969_ (.A(\adapter.game.h[4] ),
    .B(_0185_),
    .C(_0113_),
    .D(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_2 _0970_ (.A(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__or4b_1 _0971_ (.A(\adapter.game.v[8] ),
    .B(_0107_),
    .C(_0116_),
    .D_N(\adapter.game.v[9] ),
    .X(_0189_));
 sky130_fd_sc_hd__nor3_1 _0972_ (.A(_0169_),
    .B(_0115_),
    .C(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__and3_2 _0973_ (.A(net6),
    .B(_0188_),
    .C(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__and2_1 _0974_ (.A(\adapter.game.h[4] ),
    .B(_0186_),
    .X(_0192_));
 sky130_fd_sc_hd__nand3_1 _0975_ (.A(_0185_),
    .B(_0113_),
    .C(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _0976_ (.A(net6),
    .Y(_0194_));
 sky130_fd_sc_hd__or3_1 _0977_ (.A(\adapter.game.v[1] ),
    .B(\adapter.game.v[0] ),
    .C(_0116_),
    .X(_0195_));
 sky130_fd_sc_hd__or4b_1 _0978_ (.A(\adapter.game.v[8] ),
    .B(\adapter.game.v[5] ),
    .C(\adapter.game.v[4] ),
    .D_N(\adapter.game.v[9] ),
    .X(_0196_));
 sky130_fd_sc_hd__or3_1 _0979_ (.A(\adapter.game.v[7] ),
    .B(\adapter.game.v[6] ),
    .C(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or3_1 _0980_ (.A(_0194_),
    .B(_0195_),
    .C(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__nor2_1 _0981_ (.A(_0193_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__clkbuf_2 _0982_ (.A(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__buf_2 _0983_ (.A(_0078_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_2 _0984_ (.A(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__o21ai_1 _0985_ (.A1(\adapter.game.offset[0] ),
    .A2(_0200_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21oi_1 _0986_ (.A1(\adapter.game.offset[0] ),
    .A2(_0191_),
    .B1(_0203_),
    .Y(_0000_));
 sky130_fd_sc_hd__and3_1 _0987_ (.A(\adapter.game.offset[1] ),
    .B(\adapter.game.offset[0] ),
    .C(_0199_),
    .X(_0204_));
 sky130_fd_sc_hd__a21o_1 _0988_ (.A1(\adapter.game.offset[0] ),
    .A2(_0200_),
    .B1(\adapter.game.offset[1] ),
    .X(_0205_));
 sky130_fd_sc_hd__and3b_1 _0989_ (.A_N(_0204_),
    .B(_0201_),
    .C(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(_0206_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _0991_ (.A(_0145_),
    .B(_0204_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _0992_ (.A(_0145_),
    .B(_0204_),
    .Y(_0208_));
 sky130_fd_sc_hd__and3_1 _0993_ (.A(_0202_),
    .B(_0207_),
    .C(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(_0209_),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _0995_ (.A(\adapter.game.offset[3] ),
    .B(_0145_),
    .C(_0204_),
    .X(_0210_));
 sky130_fd_sc_hd__a21o_1 _0996_ (.A1(_0145_),
    .A2(_0204_),
    .B1(\adapter.game.offset[3] ),
    .X(_0211_));
 sky130_fd_sc_hd__and3b_1 _0997_ (.A_N(_0210_),
    .B(_0201_),
    .C(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(_0212_),
    .X(_0003_));
 sky130_fd_sc_hd__xnor2_1 _0999_ (.A(\adapter.game.offset[4] ),
    .B(_0210_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _1000_ (.A(net10),
    .B(_0213_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0169_),
    .B(_0188_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _1002_ (.A(_0079_),
    .B(_0190_),
    .Y(_0215_));
 sky130_fd_sc_hd__o211a_1 _1003_ (.A1(_0169_),
    .A2(_0188_),
    .B1(_0214_),
    .C1(_0215_),
    .X(_0005_));
 sky130_fd_sc_hd__and3_1 _1004_ (.A(_0094_),
    .B(\adapter.game.v[0] ),
    .C(_0187_),
    .X(_0216_));
 sky130_fd_sc_hd__or2_1 _1005_ (.A(_0079_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__a21oi_1 _1006_ (.A1(_0095_),
    .A2(_0214_),
    .B1(_0217_),
    .Y(_0006_));
 sky130_fd_sc_hd__or2_1 _1007_ (.A(_0093_),
    .B(_0216_),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_1 _1008_ (.A(_0079_),
    .B(_0188_),
    .Y(_0219_));
 sky130_fd_sc_hd__or2_1 _1009_ (.A(_0215_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _1010_ (.A(_0093_),
    .B(_0216_),
    .Y(_0221_));
 sky130_fd_sc_hd__and3_1 _1011_ (.A(_0218_),
    .B(_0220_),
    .C(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(_0222_),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _1013_ (.A(\adapter.game.v[3] ),
    .B(_0093_),
    .C(_0216_),
    .X(_0223_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(_0220_),
    .Y(_0224_));
 sky130_fd_sc_hd__a211oi_1 _1015_ (.A1(_0091_),
    .A2(_0221_),
    .B1(_0223_),
    .C1(_0224_),
    .Y(_0008_));
 sky130_fd_sc_hd__and2_1 _1016_ (.A(_0097_),
    .B(_0223_),
    .X(_0225_));
 sky130_fd_sc_hd__clkbuf_2 _1017_ (.A(_0201_),
    .X(_0226_));
 sky130_fd_sc_hd__o21ai_1 _1018_ (.A1(_0097_),
    .A2(_0223_),
    .B1(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__nor2_1 _1019_ (.A(_0225_),
    .B(_0227_),
    .Y(_0009_));
 sky130_fd_sc_hd__and3_1 _1020_ (.A(_0100_),
    .B(_0097_),
    .C(_0223_),
    .X(_0228_));
 sky130_fd_sc_hd__o21ai_1 _1021_ (.A1(_0100_),
    .A2(_0225_),
    .B1(_0226_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _1022_ (.A(_0228_),
    .B(_0229_),
    .Y(_0010_));
 sky130_fd_sc_hd__and2_1 _1023_ (.A(_0140_),
    .B(_0228_),
    .X(_0230_));
 sky130_fd_sc_hd__o21ai_1 _1024_ (.A1(_0140_),
    .A2(_0228_),
    .B1(_0226_),
    .Y(_0231_));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(_0230_),
    .B(_0231_),
    .Y(_0011_));
 sky130_fd_sc_hd__and3_1 _1026_ (.A(_0099_),
    .B(_0140_),
    .C(_0228_),
    .X(_0232_));
 sky130_fd_sc_hd__o21ai_1 _1027_ (.A1(_0099_),
    .A2(_0230_),
    .B1(_0226_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _1028_ (.A(_0232_),
    .B(_0233_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand4_1 _1029_ (.A(_0098_),
    .B(_0099_),
    .C(_0140_),
    .D(_0228_),
    .Y(_0234_));
 sky130_fd_sc_hd__buf_2 _1030_ (.A(_0202_),
    .X(_0235_));
 sky130_fd_sc_hd__o211a_1 _1031_ (.A1(_0098_),
    .A2(_0232_),
    .B1(_0234_),
    .C1(_0235_),
    .X(_0013_));
 sky130_fd_sc_hd__xor2_1 _1032_ (.A(_0090_),
    .B(_0234_),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_1 _1033_ (.A(_0224_),
    .B(_0236_),
    .Y(_0014_));
 sky130_fd_sc_hd__clkbuf_2 _1034_ (.A(\adapter.game.paddle[8] ),
    .X(_0237_));
 sky130_fd_sc_hd__xor2_1 _1035_ (.A(_0098_),
    .B(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_2 _1036_ (.A(\adapter.game.paddle[7] ),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _1037_ (.A(\adapter.game.paddle[6] ),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__a21oi_1 _1038_ (.A1(_0106_),
    .A2(_0238_),
    .B1(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__clkbuf_2 _1039_ (.A(\adapter.game.paddle[6] ),
    .X(_0242_));
 sky130_fd_sc_hd__xnor2_1 _1040_ (.A(_0099_),
    .B(_0239_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_1 _1041_ (.A(_0140_),
    .B(_0242_),
    .Y(_0244_));
 sky130_fd_sc_hd__a221o_1 _1042_ (.A1(_0242_),
    .A2(_0243_),
    .B1(_0238_),
    .B2(_0240_),
    .C1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(\adapter.game.paddle[0] ),
    .Y(_0246_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1044_ (.A(\adapter.game.paddle[5] ),
    .X(_0247_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(_0100_),
    .Y(_0248_));
 sky130_fd_sc_hd__clkbuf_2 _1046_ (.A(\adapter.game.paddle[3] ),
    .X(_0249_));
 sky130_fd_sc_hd__xor2_1 _1047_ (.A(\adapter.game.v[3] ),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a221o_1 _1048_ (.A1(_0246_),
    .A2(_0169_),
    .B1(_0247_),
    .B2(_0248_),
    .C1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_2 _1049_ (.A(\adapter.game.paddle[1] ),
    .X(_0252_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__clkbuf_2 _1051_ (.A(\adapter.game.paddle[2] ),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(_0092_),
    .Y(_0255_));
 sky130_fd_sc_hd__o22a_1 _1053_ (.A1(_0246_),
    .A2(\adapter.game.v[0] ),
    .B1(_0247_),
    .B2(_0248_),
    .X(_0256_));
 sky130_fd_sc_hd__o221a_1 _1054_ (.A1(_0094_),
    .A2(_0253_),
    .B1(_0254_),
    .B2(_0255_),
    .C1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(\adapter.game.paddle[2] ),
    .Y(_0258_));
 sky130_fd_sc_hd__clkbuf_2 _1056_ (.A(\adapter.game.paddle[4] ),
    .X(_0259_));
 sky130_fd_sc_hd__xnor2_1 _1057_ (.A(_0097_),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__o221a_1 _1058_ (.A1(_0095_),
    .A2(_0252_),
    .B1(_0258_),
    .B2(_0093_),
    .C1(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__and4bb_1 _1059_ (.A_N(_0193_),
    .B_N(_0251_),
    .C(_0257_),
    .D(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__o21ba_1 _1060_ (.A1(\adapter.game.paddle[6] ),
    .A2(_0243_),
    .B1_N(_0090_),
    .X(_0263_));
 sky130_fd_sc_hd__a31o_1 _1061_ (.A1(_0242_),
    .A2(_0239_),
    .A3(_0237_),
    .B1(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_1 _1062_ (.A(_0262_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__o31a_1 _1063_ (.A1(_0241_),
    .A2(_0245_),
    .A3(_0265_),
    .B1(\adapter.game.inPaddle ),
    .X(_0266_));
 sky130_fd_sc_hd__xnor2_1 _1064_ (.A(_0098_),
    .B(_0237_),
    .Y(_0267_));
 sky130_fd_sc_hd__and4_1 _1065_ (.A(_0262_),
    .B(_0243_),
    .C(_0267_),
    .D(_0244_),
    .X(_0268_));
 sky130_fd_sc_hd__o21a_1 _1066_ (.A1(_0266_),
    .A2(_0268_),
    .B1(_0235_),
    .X(_0015_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1067_ (.A(_0219_),
    .X(_0269_));
 sky130_fd_sc_hd__and2b_1 _1068_ (.A_N(_0170_),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _1069_ (.A(_0270_),
    .X(_0016_));
 sky130_fd_sc_hd__a21boi_1 _1070_ (.A1(_0122_),
    .A2(_0170_),
    .B1_N(_0269_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21a_1 _1071_ (.A1(_0122_),
    .A2(_0170_),
    .B1(_0271_),
    .X(_0017_));
 sky130_fd_sc_hd__and3_1 _1072_ (.A(_0122_),
    .B(_0170_),
    .C(_0120_),
    .X(_0272_));
 sky130_fd_sc_hd__a21o_1 _1073_ (.A1(_0122_),
    .A2(_0170_),
    .B1(_0120_),
    .X(_0273_));
 sky130_fd_sc_hd__and3b_1 _1074_ (.A_N(_0272_),
    .B(_0269_),
    .C(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _1075_ (.A(_0274_),
    .X(_0018_));
 sky130_fd_sc_hd__nor2_1 _1076_ (.A(_0080_),
    .B(_0186_),
    .Y(_0275_));
 sky130_fd_sc_hd__o21a_1 _1077_ (.A1(_0119_),
    .A2(_0272_),
    .B1(_0275_),
    .X(_0019_));
 sky130_fd_sc_hd__o21ai_1 _1078_ (.A1(_0083_),
    .A2(_0186_),
    .B1(_0202_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2_1 _1079_ (.A(_0192_),
    .B(_0276_),
    .Y(_0020_));
 sky130_fd_sc_hd__o21ai_1 _1080_ (.A1(_0082_),
    .A2(_0192_),
    .B1(_0269_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21oi_1 _1081_ (.A1(_0082_),
    .A2(_0192_),
    .B1(_0277_),
    .Y(_0021_));
 sky130_fd_sc_hd__and4_1 _1082_ (.A(_0082_),
    .B(_0083_),
    .C(_0084_),
    .D(_0186_),
    .X(_0278_));
 sky130_fd_sc_hd__a31o_1 _1083_ (.A1(_0082_),
    .A2(_0083_),
    .A3(_0186_),
    .B1(_0084_),
    .X(_0279_));
 sky130_fd_sc_hd__and3b_1 _1084_ (.A_N(_0278_),
    .B(_0219_),
    .C(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _1085_ (.A(_0280_),
    .X(_0022_));
 sky130_fd_sc_hd__xnor2_1 _1086_ (.A(_0081_),
    .B(_0278_),
    .Y(_0281_));
 sky130_fd_sc_hd__and2_1 _1087_ (.A(_0269_),
    .B(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _1088_ (.A(_0282_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _1089_ (.A(\adapter.game.h[7] ),
    .B(_0086_),
    .C(_0278_),
    .X(_0283_));
 sky130_fd_sc_hd__a21o_1 _1090_ (.A1(\adapter.game.h[7] ),
    .A2(_0278_),
    .B1(_0086_),
    .X(_0284_));
 sky130_fd_sc_hd__and3b_1 _1091_ (.A_N(_0283_),
    .B(_0219_),
    .C(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _1092_ (.A(_0285_),
    .X(_0024_));
 sky130_fd_sc_hd__a21boi_1 _1093_ (.A1(_0088_),
    .A2(_0283_),
    .B1_N(_0269_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21a_1 _1094_ (.A1(_0088_),
    .A2(_0283_),
    .B1(_0286_),
    .X(_0025_));
 sky130_fd_sc_hd__xnor2_1 _1095_ (.A(\adapter.game.v[3] ),
    .B(\adapter.game.ballY[2] ),
    .Y(_0287_));
 sky130_fd_sc_hd__clkbuf_2 _1096_ (.A(\adapter.game.ballY[3] ),
    .X(_0288_));
 sky130_fd_sc_hd__xnor2_1 _1097_ (.A(\adapter.game.v[4] ),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__xnor2_1 _1098_ (.A(_0099_),
    .B(\adapter.game.ballY[6] ),
    .Y(_0290_));
 sky130_fd_sc_hd__xnor2_1 _1099_ (.A(_0100_),
    .B(\adapter.game.ballY[4] ),
    .Y(_0291_));
 sky130_fd_sc_hd__and4_1 _1100_ (.A(_0287_),
    .B(_0289_),
    .C(_0290_),
    .D(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _1101_ (.A(_0092_),
    .B(\adapter.game.ballY[1] ),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _1102_ (.A(_0093_),
    .B(\adapter.game.ballY[1] ),
    .Y(_0294_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1103_ (.A(\adapter.game.ballY[0] ),
    .X(_0295_));
 sky130_fd_sc_hd__nand2_1 _1104_ (.A(_0094_),
    .B(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__or2_1 _1105_ (.A(_0094_),
    .B(_0295_),
    .X(_0297_));
 sky130_fd_sc_hd__a22o_1 _1106_ (.A1(_0293_),
    .A2(_0294_),
    .B1(_0296_),
    .B2(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__xnor2_1 _1107_ (.A(\adapter.game.v[6] ),
    .B(\adapter.game.ballY[5] ),
    .Y(_0299_));
 sky130_fd_sc_hd__xnor2_1 _1108_ (.A(_0098_),
    .B(\adapter.game.ballY[7] ),
    .Y(_0300_));
 sky130_fd_sc_hd__and3b_1 _1109_ (.A_N(_0298_),
    .B(_0299_),
    .C(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__a31o_1 _1110_ (.A1(_0188_),
    .A2(_0292_),
    .A3(_0301_),
    .B1(\adapter.game.inBallY ),
    .X(_0302_));
 sky130_fd_sc_hd__and3_1 _1111_ (.A(_0288_),
    .B(_0130_),
    .C(_0127_),
    .X(_0303_));
 sky130_fd_sc_hd__and2_1 _1112_ (.A(_0126_),
    .B(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(\adapter.game.ballY[7] ),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__o21ai_1 _1114_ (.A1(_0090_),
    .A2(_0305_),
    .B1(_0188_),
    .Y(_0306_));
 sky130_fd_sc_hd__a22o_1 _1115_ (.A1(_0128_),
    .A2(_0299_),
    .B1(_0291_),
    .B2(_0288_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_1 _1116_ (.A(\adapter.game.inBallY ),
    .B(_0287_),
    .Y(_0308_));
 sky130_fd_sc_hd__o22a_1 _1117_ (.A1(_0128_),
    .A2(_0299_),
    .B1(_0291_),
    .B2(_0288_),
    .X(_0309_));
 sky130_fd_sc_hd__or3b_1 _1118_ (.A(_0289_),
    .B(_0308_),
    .C_N(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__xnor2_1 _1119_ (.A(_0290_),
    .B(_0303_),
    .Y(_0311_));
 sky130_fd_sc_hd__or4_1 _1120_ (.A(_0298_),
    .B(_0307_),
    .C(_0310_),
    .D(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__xnor2_1 _1121_ (.A(_0300_),
    .B(_0304_),
    .Y(_0313_));
 sky130_fd_sc_hd__a2111o_1 _1122_ (.A1(_0090_),
    .A2(_0305_),
    .B1(_0306_),
    .C1(_0312_),
    .D1(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__and3_1 _1123_ (.A(_0202_),
    .B(_0302_),
    .C(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _1124_ (.A(_0315_),
    .X(_0026_));
 sky130_fd_sc_hd__buf_2 _1125_ (.A(\adapter.game.ballDirX ),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _1126_ (.A(\adapter.game.inBallX ),
    .B(_0104_),
    .Y(_0317_));
 sky130_fd_sc_hd__and3_1 _1127_ (.A(\adapter.game.inBallY ),
    .B(\adapter.game.inBallX ),
    .C(_0114_),
    .X(_0318_));
 sky130_fd_sc_hd__a211o_1 _1128_ (.A1(_0316_),
    .A2(_0317_),
    .B1(_0318_),
    .C1(_0080_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _1129_ (.A(\adapter.game.inBallY ),
    .B(_0105_),
    .Y(_0319_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1130_ (.A(\adapter.game.ballDirY ),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_2 _1131_ (.A(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _1132_ (.A1(\adapter.game.inBallY ),
    .A2(_0108_),
    .B1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__a21o_1 _1133_ (.A1(_0319_),
    .A2(_0322_),
    .B1(net10),
    .X(_0028_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1134_ (.A(\adapter.game.ballX[0] ),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_1 _1135_ (.A(_0122_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__or2_1 _1136_ (.A(\adapter.game.h[1] ),
    .B(_0323_),
    .X(_0325_));
 sky130_fd_sc_hd__xor2_1 _1137_ (.A(_0120_),
    .B(\adapter.game.ballX[1] ),
    .X(_0326_));
 sky130_fd_sc_hd__a21oi_1 _1138_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_1 _1139_ (.A(_0081_),
    .B(\adapter.game.ballX[6] ),
    .Y(_0328_));
 sky130_fd_sc_hd__and2_1 _1140_ (.A(_0081_),
    .B(\adapter.game.ballX[6] ),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_1 _1141_ (.A(_0328_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xnor2_1 _1142_ (.A(\adapter.game.h[5] ),
    .B(_0135_),
    .Y(_0331_));
 sky130_fd_sc_hd__xnor2_1 _1143_ (.A(_0084_),
    .B(\adapter.game.ballX[5] ),
    .Y(_0332_));
 sky130_fd_sc_hd__xnor2_1 _1144_ (.A(_0086_),
    .B(\adapter.game.ballX[7] ),
    .Y(_0333_));
 sky130_fd_sc_hd__and3_1 _1145_ (.A(_0331_),
    .B(_0332_),
    .C(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__xnor2_1 _1146_ (.A(_0119_),
    .B(\adapter.game.ballX[2] ),
    .Y(_0335_));
 sky130_fd_sc_hd__xnor2_1 _1147_ (.A(_0088_),
    .B(\adapter.game.ballX[8] ),
    .Y(_0336_));
 sky130_fd_sc_hd__xnor2_1 _1148_ (.A(\adapter.game.h[4] ),
    .B(_0134_),
    .Y(_0337_));
 sky130_fd_sc_hd__and3_1 _1149_ (.A(_0335_),
    .B(_0336_),
    .C(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__a41o_1 _1150_ (.A1(_0327_),
    .A2(_0330_),
    .A3(_0334_),
    .A4(_0338_),
    .B1(\adapter.game.inBallX ),
    .X(_0339_));
 sky130_fd_sc_hd__a211o_1 _1151_ (.A1(_0135_),
    .A2(_0136_),
    .B1(_0132_),
    .C1(_0133_),
    .X(_0340_));
 sky130_fd_sc_hd__a21oi_1 _1152_ (.A1(\adapter.game.ballX[8] ),
    .A2(_0340_),
    .B1(_0079_),
    .Y(_0341_));
 sky130_fd_sc_hd__and3_1 _1153_ (.A(\adapter.game.ballX[3] ),
    .B(\adapter.game.ballX[4] ),
    .C(\adapter.game.ballX[5] ),
    .X(_0342_));
 sky130_fd_sc_hd__and4_1 _1154_ (.A(_0132_),
    .B(_0133_),
    .C(_0336_),
    .D(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__o211a_1 _1155_ (.A1(_0081_),
    .A2(_0132_),
    .B1(_0333_),
    .C1(_0342_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2_1 _1156_ (.A(_0134_),
    .B(\adapter.game.ballX[4] ),
    .Y(_0345_));
 sky130_fd_sc_hd__and2_1 _1157_ (.A(_0134_),
    .B(\adapter.game.ballX[4] ),
    .X(_0346_));
 sky130_fd_sc_hd__o21ai_1 _1158_ (.A1(_0345_),
    .A2(_0346_),
    .B1(\adapter.game.h[5] ),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _1159_ (.A(_0332_),
    .Y(_0348_));
 sky130_fd_sc_hd__o32a_1 _1160_ (.A1(\adapter.game.h[5] ),
    .A2(_0345_),
    .A3(_0348_),
    .B1(_0329_),
    .B2(_0333_),
    .X(_0349_));
 sky130_fd_sc_hd__o211ai_1 _1161_ (.A1(_0330_),
    .A2(_0342_),
    .B1(_0347_),
    .C1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nor2_1 _1162_ (.A(_0332_),
    .B(_0346_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(\adapter.game.inBallX ),
    .B(_0335_),
    .Y(_0352_));
 sky130_fd_sc_hd__a31o_1 _1164_ (.A1(\adapter.game.ballX[6] ),
    .A2(_0133_),
    .A3(_0342_),
    .B1(_0336_),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _1165_ (.A(_0327_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nor4_1 _1166_ (.A(_0337_),
    .B(_0351_),
    .C(_0352_),
    .D(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__or4b_1 _1167_ (.A(_0343_),
    .B(_0344_),
    .C(_0350_),
    .D_N(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__and3_1 _1168_ (.A(_0339_),
    .B(_0341_),
    .C(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _1169_ (.A(_0357_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_2 _1170_ (.A(net2),
    .X(_0358_));
 sky130_fd_sc_hd__a21o_1 _1171_ (.A1(_0358_),
    .A2(\adapter.game.hit ),
    .B1(_0318_),
    .X(_0359_));
 sky130_fd_sc_hd__and3b_1 _1172_ (.A_N(_0268_),
    .B(_0359_),
    .C(_0201_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _1173_ (.A(_0360_),
    .X(_0030_));
 sky130_fd_sc_hd__or3b_1 _1174_ (.A(\adapter.game.v[8] ),
    .B(\adapter.game.v[0] ),
    .C_N(\adapter.game.v[9] ),
    .X(_0361_));
 sky130_fd_sc_hd__or4_1 _1175_ (.A(_0107_),
    .B(_0115_),
    .C(_0116_),
    .D(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__or3b_4 _1176_ (.A(_0194_),
    .B(_0362_),
    .C_N(_0187_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _1177_ (.A(_0358_),
    .B(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_1 _1178_ (.A(_0323_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__o211a_1 _1179_ (.A1(_0323_),
    .A2(_0200_),
    .B1(_0365_),
    .C1(_0235_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _1180_ (.A(net2),
    .B(_0363_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_2 _1181_ (.A(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(\adapter.game.ballX[1] ),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__or2_1 _1183_ (.A(_0193_),
    .B(_0198_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_2 _1184_ (.A(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_1 _1185_ (.A(\adapter.game.ballDirX ),
    .B(\adapter.game.ballX[1] ),
    .Y(_0371_));
 sky130_fd_sc_hd__or2_1 _1186_ (.A(\adapter.game.ballDirX ),
    .B(\adapter.game.ballX[1] ),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1187_ (.A1(_0371_),
    .A2(_0372_),
    .B1(_0323_),
    .Y(_0373_));
 sky130_fd_sc_hd__and3_1 _1188_ (.A(_0323_),
    .B(_0371_),
    .C(_0372_),
    .X(_0374_));
 sky130_fd_sc_hd__or3_1 _1189_ (.A(_0370_),
    .B(_0373_),
    .C(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_2 _1190_ (.A(_0080_),
    .X(_0376_));
 sky130_fd_sc_hd__a21oi_1 _1191_ (.A1(_0368_),
    .A2(_0375_),
    .B1(_0376_),
    .Y(_0032_));
 sky130_fd_sc_hd__a21boi_1 _1192_ (.A1(\adapter.game.ballX[0] ),
    .A2(_0372_),
    .B1_N(_0371_),
    .Y(_0377_));
 sky130_fd_sc_hd__xor2_1 _1193_ (.A(\adapter.game.ballDirX ),
    .B(\adapter.game.ballX[2] ),
    .X(_0378_));
 sky130_fd_sc_hd__and2_1 _1194_ (.A(_0377_),
    .B(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__nor2_1 _1195_ (.A(_0377_),
    .B(_0378_),
    .Y(_0380_));
 sky130_fd_sc_hd__or2_1 _1196_ (.A(_0379_),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_2 _1197_ (.A(_0369_),
    .X(_0382_));
 sky130_fd_sc_hd__o2bb2a_1 _1198_ (.A1_N(\adapter.game.ballX[2] ),
    .A2_N(_0367_),
    .B1(_0381_),
    .B2(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_1 _1199_ (.A(net8),
    .B(_0383_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(\adapter.game.ballDirX ),
    .Y(_0384_));
 sky130_fd_sc_hd__clkbuf_2 _1201_ (.A(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _1202_ (.A(_0385_),
    .B(_0134_),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _1203_ (.A(_0384_),
    .B(\adapter.game.ballX[3] ),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_1 _1204_ (.A(_0386_),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a21oi_1 _1205_ (.A1(_0385_),
    .A2(\adapter.game.ballX[2] ),
    .B1(_0380_),
    .Y(_0389_));
 sky130_fd_sc_hd__xnor2_1 _1206_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__o2bb2a_1 _1207_ (.A1_N(_0134_),
    .A2_N(_0367_),
    .B1(_0390_),
    .B2(_0382_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _1208_ (.A(net9),
    .B(_0391_),
    .Y(_0034_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1209_ (.A(_0366_),
    .X(_0392_));
 sky130_fd_sc_hd__o21ai_1 _1210_ (.A1(\adapter.game.ballX[2] ),
    .A2(\adapter.game.ballX[3] ),
    .B1(_0384_),
    .Y(_0393_));
 sky130_fd_sc_hd__o31a_1 _1211_ (.A1(_0377_),
    .A2(_0378_),
    .A3(_0387_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__xor2_1 _1212_ (.A(_0316_),
    .B(\adapter.game.ballX[4] ),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_1 _1213_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a21o_1 _1214_ (.A1(_0394_),
    .A2(_0395_),
    .B1(_0363_),
    .X(_0397_));
 sky130_fd_sc_hd__o2bb2a_1 _1215_ (.A1_N(_0135_),
    .A2_N(_0392_),
    .B1(_0396_),
    .B2(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_1 _1216_ (.A(net8),
    .B(_0398_),
    .Y(_0035_));
 sky130_fd_sc_hd__xor2_1 _1217_ (.A(_0316_),
    .B(_0136_),
    .X(_0399_));
 sky130_fd_sc_hd__a21o_1 _1218_ (.A1(_0385_),
    .A2(_0135_),
    .B1(_0396_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _1219_ (.A(_0399_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(_0399_),
    .B(_0400_),
    .X(_0402_));
 sky130_fd_sc_hd__nor2_1 _1221_ (.A(_0136_),
    .B(_0364_),
    .Y(_0403_));
 sky130_fd_sc_hd__a31o_1 _1222_ (.A1(_0191_),
    .A2(_0401_),
    .A3(_0402_),
    .B1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__nand2_1 _1223_ (.A(_0235_),
    .B(_0404_),
    .Y(_0036_));
 sky130_fd_sc_hd__and3_1 _1224_ (.A(_0358_),
    .B(_0132_),
    .C(_0363_),
    .X(_0405_));
 sky130_fd_sc_hd__nor3_1 _1225_ (.A(_0394_),
    .B(_0395_),
    .C(_0399_),
    .Y(_0406_));
 sky130_fd_sc_hd__o21a_1 _1226_ (.A1(_0135_),
    .A2(_0136_),
    .B1(_0385_),
    .X(_0407_));
 sky130_fd_sc_hd__xnor2_1 _1227_ (.A(_0316_),
    .B(\adapter.game.ballX[6] ),
    .Y(_0408_));
 sky130_fd_sc_hd__o21ai_1 _1228_ (.A1(_0406_),
    .A2(_0407_),
    .B1(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or3_1 _1229_ (.A(_0408_),
    .B(_0406_),
    .C(_0407_),
    .X(_0410_));
 sky130_fd_sc_hd__and3_1 _1230_ (.A(_0200_),
    .B(_0409_),
    .C(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__o21a_1 _1231_ (.A1(_0405_),
    .A2(_0411_),
    .B1(_0235_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _1232_ (.A(_0133_),
    .B(_0367_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _1233_ (.A(_0385_),
    .B(_0132_),
    .Y(_0413_));
 sky130_fd_sc_hd__xor2_1 _1234_ (.A(_0316_),
    .B(\adapter.game.ballX[7] ),
    .X(_0414_));
 sky130_fd_sc_hd__and3_1 _1235_ (.A(_0413_),
    .B(_0409_),
    .C(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a21oi_1 _1236_ (.A1(_0413_),
    .A2(_0409_),
    .B1(_0414_),
    .Y(_0416_));
 sky130_fd_sc_hd__or3_1 _1237_ (.A(_0370_),
    .B(_0415_),
    .C(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__a21oi_1 _1238_ (.A1(_0412_),
    .A2(_0417_),
    .B1(_0376_),
    .Y(_0038_));
 sky130_fd_sc_hd__buf_2 _1239_ (.A(_0080_),
    .X(_0418_));
 sky130_fd_sc_hd__inv_2 _1240_ (.A(_0414_),
    .Y(_0419_));
 sky130_fd_sc_hd__o41a_1 _1241_ (.A1(\adapter.game.ballX[4] ),
    .A2(_0136_),
    .A3(\adapter.game.ballX[6] ),
    .A4(_0133_),
    .B1(_0385_),
    .X(_0420_));
 sky130_fd_sc_hd__a31o_1 _1242_ (.A1(_0408_),
    .A2(_0406_),
    .A3(_0419_),
    .B1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__xnor2_1 _1243_ (.A(_0316_),
    .B(\adapter.game.ballX[8] ),
    .Y(_0422_));
 sky130_fd_sc_hd__xnor2_1 _1244_ (.A(_0421_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__o2bb2a_1 _1245_ (.A1_N(\adapter.game.ballX[8] ),
    .A2_N(_0392_),
    .B1(_0423_),
    .B2(_0382_),
    .X(_0424_));
 sky130_fd_sc_hd__nor2_1 _1246_ (.A(_0418_),
    .B(_0424_),
    .Y(_0039_));
 sky130_fd_sc_hd__a21oi_1 _1247_ (.A1(\adapter.game.paddle[7] ),
    .A2(_0237_),
    .B1(net3),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _1248_ (.A(net4),
    .Y(_0426_));
 sky130_fd_sc_hd__o41a_1 _1249_ (.A1(\adapter.game.paddle[5] ),
    .A2(\adapter.game.paddle[6] ),
    .A3(\adapter.game.paddle[7] ),
    .A4(\adapter.game.paddle[8] ),
    .B1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nor2_1 _1250_ (.A(_0425_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor2b_1 _1251_ (.A(_0428_),
    .B_N(_0191_),
    .Y(_0429_));
 sky130_fd_sc_hd__o211a_1 _1252_ (.A1(_0358_),
    .A2(_0429_),
    .B1(_0226_),
    .C1(\adapter.game.paddle[0] ),
    .X(_0040_));
 sky130_fd_sc_hd__or2_2 _1253_ (.A(_0363_),
    .B(_0428_),
    .X(_0430_));
 sky130_fd_sc_hd__and2_1 _1254_ (.A(net2),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_1 _1255_ (.A(_0253_),
    .B(_0430_),
    .Y(_0432_));
 sky130_fd_sc_hd__o211a_1 _1256_ (.A1(_0253_),
    .A2(_0431_),
    .B1(_0432_),
    .C1(_0235_),
    .X(_0041_));
 sky130_fd_sc_hd__o21ai_1 _1257_ (.A1(_0358_),
    .A2(_0429_),
    .B1(_0201_),
    .Y(_0433_));
 sky130_fd_sc_hd__xor2_1 _1258_ (.A(_0252_),
    .B(_0254_),
    .X(_0434_));
 sky130_fd_sc_hd__a21o_1 _1259_ (.A1(\adapter.game.paddle[7] ),
    .A2(\adapter.game.paddle[8] ),
    .B1(net3),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_2 _1260_ (.A(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_1 _1261_ (.A(_0436_),
    .B(_0427_),
    .Y(_0437_));
 sky130_fd_sc_hd__nor2_1 _1262_ (.A(_0425_),
    .B(_0434_),
    .Y(_0438_));
 sky130_fd_sc_hd__a211o_1 _1263_ (.A1(_0434_),
    .A2(_0437_),
    .B1(_0438_),
    .C1(_0363_),
    .X(_0439_));
 sky130_fd_sc_hd__o21ai_1 _1264_ (.A1(_0254_),
    .A2(_0429_),
    .B1(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _1265_ (.A(_0433_),
    .B(_0440_),
    .Y(_0042_));
 sky130_fd_sc_hd__o21ai_1 _1266_ (.A1(_0252_),
    .A2(_0254_),
    .B1(_0249_),
    .Y(_0441_));
 sky130_fd_sc_hd__or3_1 _1267_ (.A(\adapter.game.paddle[1] ),
    .B(\adapter.game.paddle[2] ),
    .C(_0249_),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _1268_ (.A(_0441_),
    .B(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__a31o_1 _1269_ (.A1(_0252_),
    .A2(_0254_),
    .A3(_0249_),
    .B1(_0436_),
    .X(_0444_));
 sky130_fd_sc_hd__a21oi_1 _1270_ (.A1(_0252_),
    .A2(_0254_),
    .B1(_0249_),
    .Y(_0445_));
 sky130_fd_sc_hd__o22a_1 _1271_ (.A1(_0437_),
    .A2(_0443_),
    .B1(_0444_),
    .B2(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__o2bb2a_1 _1272_ (.A1_N(_0249_),
    .A2_N(_0431_),
    .B1(_0446_),
    .B2(_0382_),
    .X(_0447_));
 sky130_fd_sc_hd__nor2_1 _1273_ (.A(_0418_),
    .B(_0447_),
    .Y(_0043_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(_0259_),
    .B(_0431_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _1275_ (.A(_0436_),
    .B(_0442_),
    .Y(_0449_));
 sky130_fd_sc_hd__and3_1 _1276_ (.A(_0259_),
    .B(_0444_),
    .C(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__a21oi_1 _1277_ (.A1(_0444_),
    .A2(_0449_),
    .B1(_0259_),
    .Y(_0451_));
 sky130_fd_sc_hd__or3_1 _1278_ (.A(_0430_),
    .B(_0450_),
    .C(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1279_ (.A1(_0448_),
    .A2(_0452_),
    .B1(_0376_),
    .Y(_0044_));
 sky130_fd_sc_hd__and4_1 _1280_ (.A(\adapter.game.paddle[1] ),
    .B(\adapter.game.paddle[2] ),
    .C(\adapter.game.paddle[3] ),
    .D(\adapter.game.paddle[4] ),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_1 _1281_ (.A(\adapter.game.paddle[5] ),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__or2_1 _1282_ (.A(_0247_),
    .B(_0453_),
    .X(_0455_));
 sky130_fd_sc_hd__nor3_1 _1283_ (.A(_0259_),
    .B(_0247_),
    .C(_0442_),
    .Y(_0456_));
 sky130_fd_sc_hd__o21a_1 _1284_ (.A1(_0259_),
    .A2(_0442_),
    .B1(_0247_),
    .X(_0457_));
 sky130_fd_sc_hd__o211a_1 _1285_ (.A1(_0456_),
    .A2(_0457_),
    .B1(_0436_),
    .C1(_0427_),
    .X(_0458_));
 sky130_fd_sc_hd__a31o_1 _1286_ (.A1(_0425_),
    .A2(_0454_),
    .A3(_0455_),
    .B1(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _1287_ (.A1(_0247_),
    .A2(_0431_),
    .B1(_0459_),
    .B2(_0200_),
    .X(_0460_));
 sky130_fd_sc_hd__and2_1 _1288_ (.A(_0202_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _1289_ (.A(_0461_),
    .X(_0045_));
 sky130_fd_sc_hd__or2_1 _1290_ (.A(_0435_),
    .B(_0454_),
    .X(_0462_));
 sky130_fd_sc_hd__a21bo_1 _1291_ (.A1(_0435_),
    .A2(_0456_),
    .B1_N(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__or2b_1 _1292_ (.A(_0430_),
    .B_N(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__xnor2_1 _1293_ (.A(_0242_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__or2_1 _1294_ (.A(_0433_),
    .B(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _1295_ (.A(_0466_),
    .X(_0046_));
 sky130_fd_sc_hd__a21oi_1 _1296_ (.A1(_0436_),
    .A2(_0456_),
    .B1(_0242_),
    .Y(_0467_));
 sky130_fd_sc_hd__a211oi_1 _1297_ (.A1(_0242_),
    .A2(_0462_),
    .B1(_0467_),
    .C1(_0430_),
    .Y(_0468_));
 sky130_fd_sc_hd__nor2_1 _1298_ (.A(_0239_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__a211oi_1 _1299_ (.A1(_0239_),
    .A2(_0468_),
    .B1(_0469_),
    .C1(_0433_),
    .Y(_0047_));
 sky130_fd_sc_hd__o21ai_1 _1300_ (.A1(_0358_),
    .A2(_0429_),
    .B1(_0237_),
    .Y(_0470_));
 sky130_fd_sc_hd__or3b_1 _1301_ (.A(\adapter.game.paddle[6] ),
    .B(_0239_),
    .C_N(net3),
    .X(_0471_));
 sky130_fd_sc_hd__o21a_1 _1302_ (.A1(_0240_),
    .A2(_0436_),
    .B1(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__nor2_1 _1303_ (.A(_0464_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__mux2_1 _1304_ (.A0(_0470_),
    .A1(_0237_),
    .S(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _1305_ (.A(_0418_),
    .B(_0474_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _1306_ (.A(_0295_),
    .B(_0364_),
    .Y(_0475_));
 sky130_fd_sc_hd__o211a_1 _1307_ (.A1(_0295_),
    .A2(_0200_),
    .B1(_0475_),
    .C1(_0226_),
    .X(_0049_));
 sky130_fd_sc_hd__nand2_1 _1308_ (.A(\adapter.game.ballY[1] ),
    .B(_0367_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _1309_ (.A(_0320_),
    .B(\adapter.game.ballY[1] ),
    .Y(_0477_));
 sky130_fd_sc_hd__or2_1 _1310_ (.A(\adapter.game.ballDirY ),
    .B(\adapter.game.ballY[1] ),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_1 _1311_ (.A1(_0477_),
    .A2(_0478_),
    .B1(_0295_),
    .Y(_0479_));
 sky130_fd_sc_hd__and3_1 _1312_ (.A(_0295_),
    .B(_0477_),
    .C(_0478_),
    .X(_0480_));
 sky130_fd_sc_hd__or3_1 _1313_ (.A(_0370_),
    .B(_0479_),
    .C(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a21oi_1 _1314_ (.A1(_0476_),
    .A2(_0481_),
    .B1(_0376_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand2_1 _1315_ (.A(\adapter.game.ballY[2] ),
    .B(_0367_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21bo_1 _1316_ (.A1(\adapter.game.ballY[0] ),
    .A2(_0478_),
    .B1_N(_0477_),
    .X(_0483_));
 sky130_fd_sc_hd__and2b_1 _1317_ (.A_N(\adapter.game.ballY[2] ),
    .B(\adapter.game.ballDirY ),
    .X(_0484_));
 sky130_fd_sc_hd__and2b_1 _1318_ (.A_N(_0320_),
    .B(\adapter.game.ballY[2] ),
    .X(_0485_));
 sky130_fd_sc_hd__nor2_1 _1319_ (.A(_0484_),
    .B(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__o21ai_1 _1320_ (.A1(_0483_),
    .A2(_0486_),
    .B1(_0191_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21o_1 _1321_ (.A1(_0483_),
    .A2(_0486_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__a21oi_1 _1322_ (.A1(_0482_),
    .A2(_0488_),
    .B1(_0376_),
    .Y(_0051_));
 sky130_fd_sc_hd__xor2_1 _1323_ (.A(\adapter.game.ballDirY ),
    .B(\adapter.game.ballY[3] ),
    .X(_0489_));
 sky130_fd_sc_hd__inv_2 _1324_ (.A(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__nor2_1 _1325_ (.A(_0483_),
    .B(_0485_),
    .Y(_0491_));
 sky130_fd_sc_hd__nor2_1 _1326_ (.A(_0484_),
    .B(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__xnor2_1 _1327_ (.A(_0490_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__o2bb2a_1 _1328_ (.A1_N(_0288_),
    .A2_N(_0392_),
    .B1(_0493_),
    .B2(_0382_),
    .X(_0494_));
 sky130_fd_sc_hd__nor2_1 _1329_ (.A(_0418_),
    .B(_0494_),
    .Y(_0052_));
 sky130_fd_sc_hd__o21ba_1 _1330_ (.A1(\adapter.game.ballY[2] ),
    .A2(_0288_),
    .B1_N(_0320_),
    .X(_0495_));
 sky130_fd_sc_hd__a31o_1 _1331_ (.A1(_0483_),
    .A2(_0486_),
    .A3(_0490_),
    .B1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__and2b_1 _1332_ (.A_N(_0130_),
    .B(_0320_),
    .X(_0497_));
 sky130_fd_sc_hd__and2b_1 _1333_ (.A_N(_0320_),
    .B(_0130_),
    .X(_0498_));
 sky130_fd_sc_hd__nor2_1 _1334_ (.A(_0497_),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__xnor2_1 _1335_ (.A(_0496_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o2bb2a_1 _1336_ (.A1_N(_0130_),
    .A2_N(_0392_),
    .B1(_0500_),
    .B2(_0382_),
    .X(_0501_));
 sky130_fd_sc_hd__nor2_1 _1337_ (.A(_0418_),
    .B(_0501_),
    .Y(_0053_));
 sky130_fd_sc_hd__xnor2_1 _1338_ (.A(_0321_),
    .B(_0127_),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _1339_ (.A(_0497_),
    .Y(_0503_));
 sky130_fd_sc_hd__a21oi_1 _1340_ (.A1(_0496_),
    .A2(_0503_),
    .B1(_0498_),
    .Y(_0504_));
 sky130_fd_sc_hd__xnor2_1 _1341_ (.A(_0502_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__o22a_1 _1342_ (.A1(_0127_),
    .A2(_0364_),
    .B1(_0505_),
    .B2(_0370_),
    .X(_0506_));
 sky130_fd_sc_hd__or2_1 _1343_ (.A(_0080_),
    .B(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _1344_ (.A(_0507_),
    .X(_0054_));
 sky130_fd_sc_hd__and2b_1 _1345_ (.A_N(_0321_),
    .B(_0126_),
    .X(_0508_));
 sky130_fd_sc_hd__and2b_1 _1346_ (.A_N(_0126_),
    .B(_0321_),
    .X(_0509_));
 sky130_fd_sc_hd__nor2_1 _1347_ (.A(_0508_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__o21ba_1 _1348_ (.A1(_0130_),
    .A2(_0127_),
    .B1_N(_0321_),
    .X(_0511_));
 sky130_fd_sc_hd__a31o_1 _1349_ (.A1(_0496_),
    .A2(_0499_),
    .A3(_0502_),
    .B1(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__xnor2_1 _1350_ (.A(_0510_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__o2bb2a_1 _1351_ (.A1_N(_0126_),
    .A2_N(_0392_),
    .B1(_0513_),
    .B2(_0370_),
    .X(_0514_));
 sky130_fd_sc_hd__nor2_1 _1352_ (.A(_0418_),
    .B(_0514_),
    .Y(_0055_));
 sky130_fd_sc_hd__a21o_1 _1353_ (.A1(_0510_),
    .A2(_0512_),
    .B1(_0508_),
    .X(_0515_));
 sky130_fd_sc_hd__xnor2_1 _1354_ (.A(_0321_),
    .B(\adapter.game.ballY[7] ),
    .Y(_0516_));
 sky130_fd_sc_hd__xnor2_1 _1355_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__o2bb2a_1 _1356_ (.A1_N(\adapter.game.ballY[7] ),
    .A2_N(_0392_),
    .B1(_0517_),
    .B2(_0370_),
    .X(_0518_));
 sky130_fd_sc_hd__nor2_1 _1357_ (.A(_0376_),
    .B(_0518_),
    .Y(_0056_));
 sky130_fd_sc_hd__dfxtp_1 _1358_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\adapter.game.offset[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1359_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\adapter.game.offset[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1360_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\adapter.game.offset[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1361_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\adapter.game.offset[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1362_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0004_),
    .Q(\adapter.game.offset[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1363_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0005_),
    .Q(\adapter.game.v[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1364_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\adapter.game.v[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1365_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0007_),
    .Q(\adapter.game.v[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1366_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0008_),
    .Q(\adapter.game.v[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1367_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0009_),
    .Q(\adapter.game.v[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1368_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0010_),
    .Q(\adapter.game.v[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1369_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0011_),
    .Q(\adapter.game.v[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1370_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0012_),
    .Q(\adapter.game.v[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1371_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0013_),
    .Q(\adapter.game.v[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1372_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0014_),
    .Q(\adapter.game.v[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1373_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0015_),
    .Q(\adapter.game.inPaddle ));
 sky130_fd_sc_hd__dfxtp_1 _1374_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0016_),
    .Q(\adapter.game.h[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1375_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0017_),
    .Q(\adapter.game.h[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1376_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0018_),
    .Q(\adapter.game.h[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1377_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0019_),
    .Q(\adapter.game.h[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1378_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0020_),
    .Q(\adapter.game.h[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1379_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0021_),
    .Q(\adapter.game.h[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1380_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0022_),
    .Q(\adapter.game.h[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1381_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0023_),
    .Q(\adapter.game.h[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1382_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\adapter.game.h[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1383_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0025_),
    .Q(\adapter.game.h[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1384_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0026_),
    .Q(\adapter.game.inBallY ));
 sky130_fd_sc_hd__dfxtp_1 _1385_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0027_),
    .Q(\adapter.game.ballDirX ));
 sky130_fd_sc_hd__dfxtp_1 _1386_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0028_),
    .Q(\adapter.game.ballDirY ));
 sky130_fd_sc_hd__dfxtp_1 _1387_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0029_),
    .Q(\adapter.game.inBallX ));
 sky130_fd_sc_hd__dfxtp_1 _1388_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0030_),
    .Q(\adapter.game.hit ));
 sky130_fd_sc_hd__dfxtp_1 _1389_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0031_),
    .Q(\adapter.game.ballX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1390_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0032_),
    .Q(\adapter.game.ballX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1391_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0033_),
    .Q(\adapter.game.ballX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1392_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0034_),
    .Q(\adapter.game.ballX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1393_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0035_),
    .Q(\adapter.game.ballX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1394_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0036_),
    .Q(\adapter.game.ballX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1395_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0037_),
    .Q(\adapter.game.ballX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1396_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0038_),
    .Q(\adapter.game.ballX[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1397_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0039_),
    .Q(\adapter.game.ballX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1398_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0040_),
    .Q(\adapter.game.paddle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1399_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0041_),
    .Q(\adapter.game.paddle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1400_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0042_),
    .Q(\adapter.game.paddle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1401_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0043_),
    .Q(\adapter.game.paddle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1402_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0044_),
    .Q(\adapter.game.paddle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1403_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0045_),
    .Q(\adapter.game.paddle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1404_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0046_),
    .Q(\adapter.game.paddle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1405_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0047_),
    .Q(\adapter.game.paddle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1406_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0048_),
    .Q(\adapter.game.paddle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1407_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0049_),
    .Q(\adapter.game.ballY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1408_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0050_),
    .Q(\adapter.game.ballY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1409_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0051_),
    .Q(\adapter.game.ballY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1410_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0052_),
    .Q(\adapter.game.ballY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1411_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0053_),
    .Q(\adapter.game.ballY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1412_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0054_),
    .Q(\adapter.game.ballY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1413_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0055_),
    .Q(\adapter.game.ballY[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1414_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0056_),
    .Q(\adapter.game.ballY[7] ));
 sky130_fd_sc_hd__conb_1 _1511__12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 _1512__13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 _1513__14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 _1514__15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 _1515__16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 _1516__17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 _1517__18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _1518__19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 _1519__20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 _1520__21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 _1521__22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 _1522__23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 _1523__24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 _1524__25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _1525__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _1526__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _1527__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _1528__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _1529__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _1530__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _1531__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _1532__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _1533__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _1534__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _1535__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _1536__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _1537__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _1538__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _1539__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _1540__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _1541__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _1542__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _1543__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _1544__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _1545__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _1546__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _1547__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _1548__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _1549__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _1550__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _1551__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _1552__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _1553__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _1554__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _1555__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _1564__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _1565__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _1566__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _1567__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _1568__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _1569__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _1570__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _1571__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _1572__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _1573__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _1574__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _1575__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _1576__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _1577__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _1578__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _1579__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _1580__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _1581__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _1582__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _1583__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _1584__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _1585__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _1586__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _1587__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _1588__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _1589__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _1590__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _1591__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _1592__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _1593__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _1600__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _1601__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _1602__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _1603__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _1604__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _1605__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _1606__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _1607__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _1608__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _1609__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _1610__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _1611__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _1612__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _1613__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _1614__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _1615__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _1616__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _1617__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _1618__105 (.LO(net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _1510_ (.A(net11),
    .TE_B(_0519_),
    .Z(wbs_ack_o));
 sky130_fd_sc_hd__ebufn_8 _1511_ (.A(net12),
    .TE_B(_0520_),
    .Z(wbs_dat_o[0]));
 sky130_fd_sc_hd__ebufn_8 _1512_ (.A(net13),
    .TE_B(_0521_),
    .Z(wbs_dat_o[1]));
 sky130_fd_sc_hd__ebufn_8 _1513_ (.A(net14),
    .TE_B(_0522_),
    .Z(wbs_dat_o[2]));
 sky130_fd_sc_hd__ebufn_8 _1514_ (.A(net15),
    .TE_B(_0523_),
    .Z(wbs_dat_o[3]));
 sky130_fd_sc_hd__ebufn_8 _1515_ (.A(net16),
    .TE_B(_0524_),
    .Z(wbs_dat_o[4]));
 sky130_fd_sc_hd__ebufn_8 _1516_ (.A(net17),
    .TE_B(_0525_),
    .Z(wbs_dat_o[5]));
 sky130_fd_sc_hd__ebufn_8 _1517_ (.A(net18),
    .TE_B(_0526_),
    .Z(wbs_dat_o[6]));
 sky130_fd_sc_hd__ebufn_8 _1518_ (.A(net19),
    .TE_B(_0527_),
    .Z(wbs_dat_o[7]));
 sky130_fd_sc_hd__ebufn_8 _1519_ (.A(net20),
    .TE_B(_0528_),
    .Z(wbs_dat_o[8]));
 sky130_fd_sc_hd__ebufn_8 _1520_ (.A(net21),
    .TE_B(_0529_),
    .Z(wbs_dat_o[9]));
 sky130_fd_sc_hd__ebufn_8 _1521_ (.A(net22),
    .TE_B(_0530_),
    .Z(wbs_dat_o[10]));
 sky130_fd_sc_hd__ebufn_8 _1522_ (.A(net23),
    .TE_B(_0531_),
    .Z(wbs_dat_o[11]));
 sky130_fd_sc_hd__ebufn_8 _1523_ (.A(net24),
    .TE_B(_0532_),
    .Z(wbs_dat_o[12]));
 sky130_fd_sc_hd__ebufn_8 _1524_ (.A(net25),
    .TE_B(_0533_),
    .Z(wbs_dat_o[13]));
 sky130_fd_sc_hd__ebufn_8 _1525_ (.A(net26),
    .TE_B(_0534_),
    .Z(wbs_dat_o[14]));
 sky130_fd_sc_hd__ebufn_8 _1526_ (.A(net27),
    .TE_B(_0535_),
    .Z(wbs_dat_o[15]));
 sky130_fd_sc_hd__ebufn_8 _1527_ (.A(net28),
    .TE_B(_0536_),
    .Z(wbs_dat_o[16]));
 sky130_fd_sc_hd__ebufn_8 _1528_ (.A(net29),
    .TE_B(_0537_),
    .Z(wbs_dat_o[17]));
 sky130_fd_sc_hd__ebufn_8 _1529_ (.A(net30),
    .TE_B(_0538_),
    .Z(wbs_dat_o[18]));
 sky130_fd_sc_hd__ebufn_8 _1530_ (.A(net31),
    .TE_B(_0539_),
    .Z(wbs_dat_o[19]));
 sky130_fd_sc_hd__ebufn_8 _1531_ (.A(net32),
    .TE_B(_0540_),
    .Z(wbs_dat_o[20]));
 sky130_fd_sc_hd__ebufn_8 _1532_ (.A(net33),
    .TE_B(_0541_),
    .Z(wbs_dat_o[21]));
 sky130_fd_sc_hd__ebufn_8 _1533_ (.A(net34),
    .TE_B(_0542_),
    .Z(wbs_dat_o[22]));
 sky130_fd_sc_hd__ebufn_8 _1534_ (.A(net35),
    .TE_B(_0543_),
    .Z(wbs_dat_o[23]));
 sky130_fd_sc_hd__ebufn_8 _1535_ (.A(net36),
    .TE_B(_0544_),
    .Z(wbs_dat_o[24]));
 sky130_fd_sc_hd__ebufn_8 _1536_ (.A(net37),
    .TE_B(_0545_),
    .Z(wbs_dat_o[25]));
 sky130_fd_sc_hd__ebufn_8 _1537_ (.A(net38),
    .TE_B(_0546_),
    .Z(wbs_dat_o[26]));
 sky130_fd_sc_hd__ebufn_8 _1538_ (.A(net39),
    .TE_B(_0547_),
    .Z(wbs_dat_o[27]));
 sky130_fd_sc_hd__ebufn_8 _1539_ (.A(net40),
    .TE_B(_0548_),
    .Z(wbs_dat_o[28]));
 sky130_fd_sc_hd__ebufn_8 _1540_ (.A(net41),
    .TE_B(_0549_),
    .Z(wbs_dat_o[29]));
 sky130_fd_sc_hd__ebufn_8 _1541_ (.A(net42),
    .TE_B(_0550_),
    .Z(wbs_dat_o[30]));
 sky130_fd_sc_hd__ebufn_8 _1542_ (.A(net43),
    .TE_B(_0551_),
    .Z(wbs_dat_o[31]));
 sky130_fd_sc_hd__ebufn_8 _1543_ (.A(net44),
    .TE_B(_0552_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1544_ (.A(net45),
    .TE_B(_0553_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1545_ (.A(net46),
    .TE_B(_0554_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1546_ (.A(net47),
    .TE_B(_0555_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1547_ (.A(net48),
    .TE_B(_0556_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1548_ (.A(net49),
    .TE_B(_0557_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1549_ (.A(net50),
    .TE_B(_0558_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1550_ (.A(net51),
    .TE_B(_0559_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1551_ (.A(net52),
    .TE_B(_0560_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1552_ (.A(net53),
    .TE_B(_0561_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1553_ (.A(net54),
    .TE_B(_0562_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1554_ (.A(net55),
    .TE_B(_0563_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1555_ (.A(net56),
    .TE_B(_0564_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1556_ (.A(\adapter.game.red ),
    .TE_B(_0565_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1557_ (.A(\adapter.game.green ),
    .TE_B(_0566_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1558_ (.A(\adapter.blue ),
    .TE_B(_0567_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1559_ (.A(\adapter.game.hsync ),
    .TE_B(_0568_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1560_ (.A(\adapter.game.vsync ),
    .TE_B(_0569_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1561_ (.A(\adapter.game.speaker ),
    .TE_B(_0570_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1562_ (.A(net8),
    .TE_B(_0571_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1563_ (.A(net1),
    .TE_B(_0572_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1564_ (.A(net57),
    .TE_B(_0573_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1565_ (.A(net58),
    .TE_B(_0574_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1566_ (.A(net59),
    .TE_B(_0575_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1567_ (.A(net60),
    .TE_B(_0576_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1568_ (.A(net61),
    .TE_B(_0577_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1569_ (.A(net62),
    .TE_B(_0578_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1570_ (.A(net63),
    .TE_B(_0579_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1571_ (.A(net64),
    .TE_B(_0580_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1572_ (.A(net65),
    .TE_B(_0581_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1573_ (.A(net66),
    .TE_B(_0582_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1574_ (.A(net67),
    .TE_B(_0583_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1575_ (.A(net68),
    .TE_B(_0584_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _1576_ (.A(net69),
    .TE_B(_0585_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _1577_ (.A(net70),
    .TE_B(_0586_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _1578_ (.A(net71),
    .TE_B(_0587_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _1579_ (.A(net72),
    .TE_B(_0588_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _1580_ (.A(net73),
    .TE_B(_0589_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _1581_ (.A(net74),
    .TE_B(_0590_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _1582_ (.A(net75),
    .TE_B(_0591_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _1583_ (.A(net76),
    .TE_B(_0592_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _1584_ (.A(net77),
    .TE_B(_0593_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _1585_ (.A(net78),
    .TE_B(_0594_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _1586_ (.A(net79),
    .TE_B(_0595_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _1587_ (.A(net80),
    .TE_B(_0596_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _1588_ (.A(net81),
    .TE_B(_0597_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _1589_ (.A(net82),
    .TE_B(_0598_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _1590_ (.A(net83),
    .TE_B(_0599_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _1591_ (.A(net84),
    .TE_B(_0600_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _1592_ (.A(net85),
    .TE_B(_0601_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _1593_ (.A(net86),
    .TE_B(_0602_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _1594_ (.A(net8),
    .TE_B(_0603_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _1595_ (.A(net8),
    .TE_B(_0604_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _1596_ (.A(net9),
    .TE_B(_0605_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _1597_ (.A(net10),
    .TE_B(_0606_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _1598_ (.A(net10),
    .TE_B(_0607_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _1599_ (.A(net8),
    .TE_B(_0608_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _1600_ (.A(net87),
    .TE_B(_0609_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _1601_ (.A(net88),
    .TE_B(_0610_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _1602_ (.A(net89),
    .TE_B(_0611_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _1603_ (.A(net90),
    .TE_B(_0612_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _1604_ (.A(net91),
    .TE_B(_0613_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _1605_ (.A(net92),
    .TE_B(_0614_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _1606_ (.A(net93),
    .TE_B(_0615_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _1607_ (.A(net94),
    .TE_B(_0616_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _1608_ (.A(net95),
    .TE_B(_0617_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _1609_ (.A(net96),
    .TE_B(_0618_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _1610_ (.A(net97),
    .TE_B(_0619_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _1611_ (.A(net98),
    .TE_B(_0620_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _1612_ (.A(net99),
    .TE_B(_0621_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _1613_ (.A(net100),
    .TE_B(_0622_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _1614_ (.A(net101),
    .TE_B(_0623_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _1615_ (.A(net102),
    .TE_B(_0624_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _1616_ (.A(net103),
    .TE_B(_0625_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _1617_ (.A(net104),
    .TE_B(_0626_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _1618_ (.A(net105),
    .TE_B(_0627_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(io_in[8]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[9]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(wb_rst_i),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(\adapter.debug_design_reset ),
    .X(net10));
 sky130_fd_sc_hd__conb_1 _1510__11 (.LO(net11));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
endmodule

