magic
tech sky130A
magscale 1 2
timestamp 1680612644
<< viali >>
rect 1869 37281 1903 37315
rect 18245 37281 18279 37315
rect 25789 37281 25823 37315
rect 28641 37281 28675 37315
rect 30389 37281 30423 37315
rect 32965 37281 32999 37315
rect 38301 37281 38335 37315
rect 1685 37213 1719 37247
rect 2513 37213 2547 37247
rect 3433 37213 3467 37247
rect 4169 37213 4203 37247
rect 4813 37213 4847 37247
rect 6561 37213 6595 37247
rect 9229 37213 9263 37247
rect 14473 37213 14507 37247
rect 14933 37213 14967 37247
rect 15761 37213 15795 37247
rect 17601 37213 17635 37247
rect 18889 37213 18923 37247
rect 19809 37213 19843 37247
rect 21005 37213 21039 37247
rect 22109 37213 22143 37247
rect 22753 37213 22787 37247
rect 23581 37213 23615 37247
rect 26617 37213 26651 37247
rect 27169 37213 27203 37247
rect 27813 37213 27847 37247
rect 29929 37213 29963 37247
rect 32505 37213 32539 37247
rect 36921 37213 36955 37247
rect 38025 37213 38059 37247
rect 26433 37145 26467 37179
rect 30113 37145 30147 37179
rect 32689 37145 32723 37179
rect 35081 37145 35115 37179
rect 36737 37145 36771 37179
rect 4721 37077 4755 37111
rect 15669 37077 15703 37111
rect 17509 37077 17543 37111
rect 22201 37077 22235 37111
rect 38209 36873 38243 36907
rect 1869 36805 1903 36839
rect 4353 36805 4387 36839
rect 14657 36805 14691 36839
rect 16313 36805 16347 36839
rect 22293 36805 22327 36839
rect 32505 36805 32539 36839
rect 3709 36737 3743 36771
rect 4169 36737 4203 36771
rect 6561 36737 6595 36771
rect 9229 36737 9263 36771
rect 19165 36737 19199 36771
rect 19625 36737 19659 36771
rect 24409 36737 24443 36771
rect 27169 36737 27203 36771
rect 38117 36737 38151 36771
rect 3525 36669 3559 36703
rect 4629 36669 4663 36703
rect 6745 36669 6779 36703
rect 7113 36669 7147 36703
rect 9413 36669 9447 36703
rect 9689 36669 9723 36703
rect 14473 36669 14507 36703
rect 18061 36669 18095 36703
rect 18981 36669 19015 36703
rect 19809 36669 19843 36703
rect 20729 36669 20763 36703
rect 22109 36669 22143 36703
rect 22845 36669 22879 36703
rect 24593 36669 24627 36703
rect 24869 36669 24903 36703
rect 27353 36669 27387 36703
rect 27629 36669 27663 36703
rect 29469 36669 29503 36703
rect 29653 36669 29687 36703
rect 29929 36669 29963 36703
rect 32321 36669 32355 36703
rect 32781 36669 32815 36703
rect 34621 36669 34655 36703
rect 34805 36669 34839 36703
rect 35081 36669 35115 36703
rect 37473 36533 37507 36567
rect 6469 36329 6503 36363
rect 9413 36329 9447 36363
rect 19901 36329 19935 36363
rect 23397 36329 23431 36363
rect 2789 36193 2823 36227
rect 3985 36193 4019 36227
rect 4445 36193 4479 36227
rect 14749 36193 14783 36227
rect 16129 36193 16163 36227
rect 17417 36193 17451 36227
rect 18705 36193 18739 36227
rect 18889 36193 18923 36227
rect 21005 36193 21039 36227
rect 22109 36193 22143 36227
rect 25145 36193 25179 36227
rect 27353 36193 27387 36227
rect 30205 36193 30239 36227
rect 32505 36193 32539 36227
rect 36737 36193 36771 36227
rect 37197 36193 37231 36227
rect 1593 36125 1627 36159
rect 6377 36125 6411 36159
rect 9321 36125 9355 36159
rect 19993 36125 20027 36159
rect 23305 36125 23339 36159
rect 24593 36125 24627 36159
rect 26893 36125 26927 36159
rect 29745 36125 29779 36159
rect 32045 36125 32079 36159
rect 37657 36125 37691 36159
rect 1777 36057 1811 36091
rect 4169 36057 4203 36091
rect 14933 36057 14967 36091
rect 21189 36057 21223 36091
rect 24777 36057 24811 36091
rect 27077 36057 27111 36091
rect 29929 36057 29963 36091
rect 32229 36057 32263 36091
rect 37013 36057 37047 36091
rect 37749 36057 37783 36091
rect 2421 35785 2455 35819
rect 3065 35785 3099 35819
rect 3709 35785 3743 35819
rect 15117 35785 15151 35819
rect 18797 35785 18831 35819
rect 21097 35785 21131 35819
rect 23673 35785 23707 35819
rect 25145 35785 25179 35819
rect 30021 35785 30055 35819
rect 30665 35785 30699 35819
rect 26065 35717 26099 35751
rect 27629 35717 27663 35751
rect 34437 35717 34471 35751
rect 1685 35649 1719 35683
rect 2513 35649 2547 35683
rect 3157 35649 3191 35683
rect 3617 35649 3651 35683
rect 15209 35649 15243 35683
rect 17121 35649 17155 35683
rect 18889 35649 18923 35683
rect 21005 35649 21039 35683
rect 23581 35649 23615 35683
rect 24409 35649 24443 35683
rect 25053 35649 25087 35683
rect 25973 35649 26007 35683
rect 29469 35649 29503 35683
rect 30113 35649 30147 35683
rect 30573 35649 30607 35683
rect 31401 35649 31435 35683
rect 38117 35649 38151 35683
rect 16865 35581 16899 35615
rect 29285 35581 29319 35615
rect 33057 35581 33091 35615
rect 34621 35581 34655 35615
rect 35725 35581 35759 35615
rect 36737 35581 36771 35615
rect 36921 35581 36955 35615
rect 37473 35581 37507 35615
rect 18245 35445 18279 35479
rect 38209 35445 38243 35479
rect 16957 35241 16991 35275
rect 18705 35241 18739 35275
rect 26617 35241 26651 35275
rect 27169 35241 27203 35275
rect 27997 35241 28031 35275
rect 28641 35241 28675 35275
rect 30113 35241 30147 35275
rect 30665 35241 30699 35275
rect 31769 35241 31803 35275
rect 32321 35241 32355 35275
rect 33057 35241 33091 35275
rect 34345 35241 34379 35275
rect 34989 35241 35023 35275
rect 35725 35241 35759 35275
rect 19533 35105 19567 35139
rect 37841 35105 37875 35139
rect 14289 35037 14323 35071
rect 17141 35037 17175 35071
rect 19625 35037 19659 35071
rect 20637 35037 20671 35071
rect 21281 35037 21315 35071
rect 26525 35037 26559 35071
rect 28089 35037 28123 35071
rect 28549 35037 28583 35071
rect 30021 35037 30055 35071
rect 31677 35037 31711 35071
rect 33149 35037 33183 35071
rect 35081 35037 35115 35071
rect 35633 35037 35667 35071
rect 38301 35037 38335 35071
rect 14556 34969 14590 35003
rect 18689 34969 18723 35003
rect 18889 34969 18923 35003
rect 21526 34969 21560 35003
rect 38117 34969 38151 35003
rect 15669 34901 15703 34935
rect 18521 34901 18555 34935
rect 19993 34901 20027 34935
rect 20821 34901 20855 34935
rect 22661 34901 22695 34935
rect 17601 34697 17635 34731
rect 21005 34697 21039 34731
rect 37565 34697 37599 34731
rect 17785 34629 17819 34663
rect 36737 34629 36771 34663
rect 2513 34561 2547 34595
rect 18153 34561 18187 34595
rect 18705 34561 18739 34595
rect 20821 34561 20855 34595
rect 22937 34561 22971 34595
rect 33701 34561 33735 34595
rect 37473 34561 37507 34595
rect 38301 34561 38335 34595
rect 3341 34493 3375 34527
rect 14933 34493 14967 34527
rect 19901 34493 19935 34527
rect 20177 34493 20211 34527
rect 20637 34493 20671 34527
rect 23029 34493 23063 34527
rect 23581 34493 23615 34527
rect 23765 34493 23799 34527
rect 24501 34493 24535 34527
rect 35725 34493 35759 34527
rect 36921 34493 36955 34527
rect 14657 34425 14691 34459
rect 28457 34425 28491 34459
rect 29101 34425 29135 34459
rect 32689 34425 32723 34459
rect 14473 34357 14507 34391
rect 17785 34357 17819 34391
rect 18797 34357 18831 34391
rect 33793 34357 33827 34391
rect 14657 34153 14691 34187
rect 17049 34153 17083 34187
rect 18429 34153 18463 34187
rect 20361 34153 20395 34187
rect 23397 34153 23431 34187
rect 35173 34153 35207 34187
rect 36001 34153 36035 34187
rect 15117 34017 15151 34051
rect 26985 34017 27019 34051
rect 32229 34017 32263 34051
rect 34069 34017 34103 34051
rect 38301 34017 38335 34051
rect 1961 33949 1995 33983
rect 2789 33949 2823 33983
rect 14473 33949 14507 33983
rect 15393 33949 15427 33983
rect 16865 33949 16899 33983
rect 17141 33949 17175 33983
rect 18613 33949 18647 33983
rect 18889 33949 18923 33983
rect 19993 33949 20027 33983
rect 21465 33949 21499 33983
rect 23305 33949 23339 33983
rect 25973 33949 26007 33983
rect 27169 33949 27203 33983
rect 27813 33949 27847 33983
rect 27997 33949 28031 33983
rect 36461 33949 36495 33983
rect 20361 33881 20395 33915
rect 21710 33881 21744 33915
rect 25706 33881 25740 33915
rect 27353 33881 27387 33915
rect 32413 33881 32447 33915
rect 36645 33881 36679 33915
rect 2697 33813 2731 33847
rect 16681 33813 16715 33847
rect 18797 33813 18831 33847
rect 20545 33813 20579 33847
rect 22845 33813 22879 33847
rect 24593 33813 24627 33847
rect 27905 33813 27939 33847
rect 17141 33609 17175 33643
rect 19717 33609 19751 33643
rect 21281 33609 21315 33643
rect 23765 33609 23799 33643
rect 25513 33609 25547 33643
rect 27261 33609 27295 33643
rect 32413 33609 32447 33643
rect 36185 33609 36219 33643
rect 36829 33609 36863 33643
rect 2053 33541 2087 33575
rect 17233 33541 17267 33575
rect 24501 33541 24535 33575
rect 24717 33541 24751 33575
rect 33793 33541 33827 33575
rect 1869 33473 1903 33507
rect 15025 33473 15059 33507
rect 15117 33473 15151 33507
rect 17325 33473 17359 33507
rect 19901 33473 19935 33507
rect 19993 33473 20027 33507
rect 20085 33473 20119 33507
rect 21097 33473 21131 33507
rect 23673 33473 23707 33507
rect 25329 33473 25363 33507
rect 27169 33473 27203 33507
rect 27353 33473 27387 33507
rect 27905 33473 27939 33507
rect 32321 33473 32355 33507
rect 36277 33473 36311 33507
rect 36921 33473 36955 33507
rect 38117 33473 38151 33507
rect 2789 33405 2823 33439
rect 14657 33405 14691 33439
rect 16865 33405 16899 33439
rect 33609 33405 33643 33439
rect 34529 33405 34563 33439
rect 20269 33337 20303 33371
rect 24869 33337 24903 33371
rect 14841 33269 14875 33303
rect 24685 33269 24719 33303
rect 27997 33269 28031 33303
rect 37473 33269 37507 33303
rect 21005 33065 21039 33099
rect 26157 33065 26191 33099
rect 26801 33065 26835 33099
rect 24869 32997 24903 33031
rect 26341 32997 26375 33031
rect 20258 32929 20292 32963
rect 21281 32929 21315 32963
rect 21465 32929 21499 32963
rect 22293 32929 22327 32963
rect 24961 32929 24995 32963
rect 28181 32929 28215 32963
rect 36461 32929 36495 32963
rect 38301 32929 38335 32963
rect 2237 32861 2271 32895
rect 10425 32861 10459 32895
rect 10609 32861 10643 32895
rect 12909 32861 12943 32895
rect 14381 32861 14415 32895
rect 16313 32861 16347 32895
rect 18245 32861 18279 32895
rect 20178 32861 20212 32895
rect 20361 32861 20395 32895
rect 20453 32861 20487 32895
rect 21189 32861 21223 32895
rect 21373 32861 21407 32895
rect 22385 32861 22419 32895
rect 22937 32861 22971 32895
rect 23121 32861 23155 32895
rect 26065 32861 26099 32895
rect 26157 32861 26191 32895
rect 27077 32861 27111 32895
rect 27169 32861 27203 32895
rect 27261 32861 27295 32895
rect 27445 32861 27479 32895
rect 27905 32861 27939 32895
rect 28089 32861 28123 32895
rect 28273 32861 28307 32895
rect 28365 32861 28399 32895
rect 14648 32793 14682 32827
rect 16580 32793 16614 32827
rect 18429 32793 18463 32827
rect 22109 32793 22143 32827
rect 24777 32793 24811 32827
rect 25145 32793 25179 32827
rect 25697 32793 25731 32827
rect 36645 32793 36679 32827
rect 10517 32725 10551 32759
rect 12725 32725 12759 32759
rect 15761 32725 15795 32759
rect 17693 32725 17727 32759
rect 19993 32725 20027 32759
rect 22385 32725 22419 32759
rect 25053 32725 25087 32759
rect 28549 32725 28583 32759
rect 14657 32521 14691 32555
rect 24685 32521 24719 32555
rect 27537 32521 27571 32555
rect 36553 32521 36587 32555
rect 3893 32385 3927 32419
rect 10894 32385 10928 32419
rect 12440 32385 12474 32419
rect 14841 32385 14875 32419
rect 15117 32385 15151 32419
rect 17417 32385 17451 32419
rect 17601 32385 17635 32419
rect 18245 32385 18279 32419
rect 18521 32385 18555 32419
rect 19441 32385 19475 32419
rect 19901 32385 19935 32419
rect 24869 32385 24903 32419
rect 25099 32385 25133 32419
rect 27169 32385 27203 32419
rect 27261 32385 27295 32419
rect 27537 32385 27571 32419
rect 29009 32385 29043 32419
rect 36461 32385 36495 32419
rect 37657 32385 37691 32419
rect 2697 32317 2731 32351
rect 3709 32317 3743 32351
rect 8677 32317 8711 32351
rect 11161 32317 11195 32351
rect 12173 32317 12207 32351
rect 18061 32317 18095 32351
rect 19625 32317 19659 32351
rect 21189 32317 21223 32351
rect 21465 32317 21499 32351
rect 24961 32317 24995 32351
rect 25237 32317 25271 32351
rect 25329 32317 25363 32351
rect 27445 32317 27479 32351
rect 29101 32317 29135 32351
rect 9045 32249 9079 32283
rect 9781 32249 9815 32283
rect 19257 32249 19291 32283
rect 28641 32249 28675 32283
rect 9137 32181 9171 32215
rect 13553 32181 13587 32215
rect 15025 32181 15059 32215
rect 17233 32181 17267 32215
rect 18429 32181 18463 32215
rect 19625 32181 19659 32215
rect 10425 31977 10459 32011
rect 19625 31977 19659 32011
rect 24777 31977 24811 32011
rect 24961 31977 24995 32011
rect 27077 31977 27111 32011
rect 27905 31977 27939 32011
rect 28549 31977 28583 32011
rect 31125 31977 31159 32011
rect 4445 31909 4479 31943
rect 15025 31909 15059 31943
rect 18153 31909 18187 31943
rect 22845 31909 22879 31943
rect 27721 31909 27755 31943
rect 10241 31841 10275 31875
rect 13553 31841 13587 31875
rect 16957 31841 16991 31875
rect 20545 31841 20579 31875
rect 20637 31841 20671 31875
rect 20913 31841 20947 31875
rect 21465 31841 21499 31875
rect 23581 31841 23615 31875
rect 26985 31841 27019 31875
rect 27169 31841 27203 31875
rect 1685 31773 1719 31807
rect 2513 31773 2547 31807
rect 4629 31773 4663 31807
rect 10149 31773 10183 31807
rect 13297 31773 13331 31807
rect 15393 31773 15427 31807
rect 15577 31773 15611 31807
rect 16773 31773 16807 31807
rect 18429 31773 18463 31807
rect 19533 31773 19567 31807
rect 19717 31773 19751 31807
rect 19809 31773 19843 31807
rect 20453 31773 20487 31807
rect 20729 31773 20763 31807
rect 21721 31773 21755 31807
rect 23489 31773 23523 31807
rect 27261 31773 27295 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 29745 31773 29779 31807
rect 33793 31773 33827 31807
rect 9413 31705 9447 31739
rect 15301 31705 15335 31739
rect 18153 31705 18187 31739
rect 24593 31705 24627 31739
rect 27873 31705 27907 31739
rect 28089 31705 28123 31739
rect 30012 31705 30046 31739
rect 2421 31637 2455 31671
rect 9321 31637 9355 31671
rect 12173 31637 12207 31671
rect 15209 31637 15243 31671
rect 18337 31637 18371 31671
rect 23857 31637 23891 31671
rect 24793 31637 24827 31671
rect 33885 31637 33919 31671
rect 3525 31433 3559 31467
rect 14657 31433 14691 31467
rect 18153 31433 18187 31467
rect 24593 31433 24627 31467
rect 25145 31433 25179 31467
rect 26249 31433 26283 31467
rect 27813 31433 27847 31467
rect 30113 31433 30147 31467
rect 14841 31365 14875 31399
rect 15669 31365 15703 31399
rect 25973 31365 26007 31399
rect 34069 31365 34103 31399
rect 35725 31365 35759 31399
rect 2329 31297 2363 31331
rect 3617 31297 3651 31331
rect 9505 31297 9539 31331
rect 9689 31297 9723 31331
rect 15853 31297 15887 31331
rect 16037 31297 16071 31331
rect 16129 31297 16163 31331
rect 18429 31297 18463 31331
rect 24409 31297 24443 31331
rect 24593 31297 24627 31331
rect 25053 31297 25087 31331
rect 25237 31297 25271 31331
rect 25881 31297 25915 31331
rect 26065 31297 26099 31331
rect 27445 31297 27479 31331
rect 30021 31297 30055 31331
rect 30205 31297 30239 31331
rect 8585 31229 8619 31263
rect 18153 31229 18187 31263
rect 18337 31229 18371 31263
rect 27537 31229 27571 31263
rect 33885 31229 33919 31263
rect 2237 31161 2271 31195
rect 8953 31161 8987 31195
rect 15209 31161 15243 31195
rect 25697 31161 25731 31195
rect 2973 31093 3007 31127
rect 4077 31093 4111 31127
rect 9045 31093 9079 31127
rect 9505 31093 9539 31127
rect 14841 31093 14875 31127
rect 37841 31093 37875 31127
rect 4537 30889 4571 30923
rect 14289 30889 14323 30923
rect 22385 30889 22419 30923
rect 25605 30889 25639 30923
rect 27813 30889 27847 30923
rect 30113 30889 30147 30923
rect 13553 30821 13587 30855
rect 14657 30821 14691 30855
rect 1593 30753 1627 30787
rect 1777 30753 1811 30787
rect 2789 30753 2823 30787
rect 13737 30753 13771 30787
rect 14749 30753 14783 30787
rect 15669 30753 15703 30787
rect 19441 30753 19475 30787
rect 19625 30753 19659 30787
rect 25881 30753 25915 30787
rect 26065 30753 26099 30787
rect 37841 30753 37875 30787
rect 38301 30753 38335 30787
rect 10793 30685 10827 30719
rect 11069 30685 11103 30719
rect 13461 30685 13495 30719
rect 14473 30685 14507 30719
rect 17877 30685 17911 30719
rect 17969 30685 18003 30719
rect 18153 30685 18187 30719
rect 18613 30685 18647 30719
rect 18797 30685 18831 30719
rect 19717 30685 19751 30719
rect 22109 30685 22143 30719
rect 25789 30685 25823 30719
rect 25973 30685 26007 30719
rect 27629 30685 27663 30719
rect 27813 30685 27847 30719
rect 4445 30617 4479 30651
rect 17417 30617 17451 30651
rect 19441 30617 19475 30651
rect 22385 30617 22419 30651
rect 30021 30617 30055 30651
rect 38117 30617 38151 30651
rect 13737 30549 13771 30583
rect 18061 30549 18095 30583
rect 18705 30549 18739 30583
rect 22201 30549 22235 30583
rect 15209 30345 15243 30379
rect 15377 30345 15411 30379
rect 17325 30345 17359 30379
rect 37657 30345 37691 30379
rect 15577 30277 15611 30311
rect 17141 30277 17175 30311
rect 17233 30277 17267 30311
rect 18337 30277 18371 30311
rect 19441 30277 19475 30311
rect 19533 30277 19567 30311
rect 23121 30277 23155 30311
rect 30639 30277 30673 30311
rect 2973 30209 3007 30243
rect 4077 30209 4111 30243
rect 8125 30209 8159 30243
rect 8769 30209 8803 30243
rect 10149 30209 10183 30243
rect 11897 30209 11931 30243
rect 12081 30209 12115 30243
rect 12173 30209 12207 30243
rect 14565 30209 14599 30243
rect 18153 30209 18187 30243
rect 19625 30209 19659 30243
rect 20545 30209 20579 30243
rect 22385 30209 22419 30243
rect 23029 30209 23063 30243
rect 23213 30209 23247 30243
rect 23857 30209 23891 30243
rect 25973 30209 26007 30243
rect 27721 30209 27755 30243
rect 27905 30209 27939 30243
rect 29673 30209 29707 30243
rect 29929 30209 29963 30243
rect 30514 30209 30548 30243
rect 31493 30209 31527 30243
rect 31585 30209 31619 30243
rect 31769 30209 31803 30243
rect 32689 30209 32723 30243
rect 37565 30209 37599 30243
rect 4261 30141 4295 30175
rect 4721 30141 4755 30175
rect 8861 30141 8895 30175
rect 10701 30141 10735 30175
rect 13185 30141 13219 30175
rect 17969 30141 18003 30175
rect 20269 30141 20303 30175
rect 22477 30141 22511 30175
rect 23949 30141 23983 30175
rect 26065 30141 26099 30175
rect 28089 30141 28123 30175
rect 31033 30141 31067 30175
rect 32597 30141 32631 30175
rect 9137 30073 9171 30107
rect 13553 30073 13587 30107
rect 14749 30073 14783 30107
rect 17509 30073 17543 30107
rect 19257 30073 19291 30107
rect 22017 30073 22051 30107
rect 24225 30073 24259 30107
rect 26341 30073 26375 30107
rect 31769 30073 31803 30107
rect 2145 30005 2179 30039
rect 2881 30005 2915 30039
rect 7665 30005 7699 30039
rect 8033 30005 8067 30039
rect 11713 30005 11747 30039
rect 13645 30005 13679 30039
rect 15393 30005 15427 30039
rect 16957 30005 16991 30039
rect 19809 30005 19843 30039
rect 28549 30005 28583 30039
rect 30389 30005 30423 30039
rect 30941 30005 30975 30039
rect 32413 30005 32447 30039
rect 4445 29801 4479 29835
rect 5365 29801 5399 29835
rect 12081 29801 12115 29835
rect 19809 29801 19843 29835
rect 20637 29801 20671 29835
rect 21833 29801 21867 29835
rect 25053 29801 25087 29835
rect 28457 29801 28491 29835
rect 28641 29801 28675 29835
rect 29929 29801 29963 29835
rect 30573 29801 30607 29835
rect 9137 29733 9171 29767
rect 14289 29733 14323 29767
rect 17877 29733 17911 29767
rect 3433 29665 3467 29699
rect 19625 29665 19659 29699
rect 24685 29665 24719 29699
rect 26709 29665 26743 29699
rect 31125 29665 31159 29699
rect 37197 29665 37231 29699
rect 4537 29597 4571 29631
rect 9321 29597 9355 29631
rect 9413 29597 9447 29631
rect 10057 29597 10091 29631
rect 10701 29597 10735 29631
rect 12541 29597 12575 29631
rect 13461 29597 13495 29631
rect 13737 29597 13771 29631
rect 14448 29597 14482 29631
rect 14785 29597 14819 29631
rect 14933 29597 14967 29631
rect 15577 29597 15611 29631
rect 15761 29597 15795 29631
rect 17417 29597 17451 29631
rect 19717 29597 19751 29631
rect 19993 29597 20027 29631
rect 20637 29597 20671 29631
rect 20821 29597 20855 29631
rect 24777 29597 24811 29631
rect 26525 29597 26559 29631
rect 29745 29597 29779 29631
rect 29929 29597 29963 29631
rect 30754 29597 30788 29631
rect 31217 29597 31251 29631
rect 32137 29597 32171 29631
rect 38301 29597 38335 29631
rect 1593 29529 1627 29563
rect 3249 29529 3283 29563
rect 5089 29529 5123 29563
rect 9137 29529 9171 29563
rect 10946 29529 10980 29563
rect 14565 29529 14599 29563
rect 14657 29529 14691 29563
rect 17325 29529 17359 29563
rect 17877 29529 17911 29563
rect 22017 29529 22051 29563
rect 22201 29529 22235 29563
rect 27261 29529 27295 29563
rect 28825 29529 28859 29563
rect 32321 29529 32355 29563
rect 32505 29529 32539 29563
rect 38117 29529 38151 29563
rect 10241 29461 10275 29495
rect 12633 29461 12667 29495
rect 13277 29461 13311 29495
rect 13645 29461 13679 29495
rect 15393 29461 15427 29495
rect 17141 29461 17175 29495
rect 19901 29461 19935 29495
rect 27353 29461 27387 29495
rect 28625 29461 28659 29495
rect 30757 29461 30791 29495
rect 11713 29257 11747 29291
rect 11897 29257 11931 29291
rect 31585 29257 31619 29291
rect 18328 29189 18362 29223
rect 25145 29189 25179 29223
rect 30757 29189 30791 29223
rect 31401 29189 31435 29223
rect 2145 29121 2179 29155
rect 4813 29121 4847 29155
rect 8217 29121 8251 29155
rect 10425 29121 10459 29155
rect 10977 29121 11011 29155
rect 12265 29121 12299 29155
rect 13369 29121 13403 29155
rect 15025 29121 15059 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 21005 29121 21039 29155
rect 21189 29121 21223 29155
rect 23397 29121 23431 29155
rect 26433 29121 26467 29155
rect 30573 29121 30607 29155
rect 31217 29121 31251 29155
rect 37841 29121 37875 29155
rect 2329 29053 2363 29087
rect 2881 29053 2915 29087
rect 8125 29053 8159 29087
rect 13829 29053 13863 29087
rect 14565 29053 14599 29087
rect 15945 29053 15979 29087
rect 18061 29053 18095 29087
rect 30389 29053 30423 29087
rect 15485 28985 15519 29019
rect 15577 28985 15611 29019
rect 16865 28985 16899 29019
rect 19441 28985 19475 29019
rect 26249 28985 26283 29019
rect 4721 28917 4755 28951
rect 7849 28917 7883 28951
rect 11897 28917 11931 28951
rect 13645 28917 13679 28951
rect 14933 28917 14967 28951
rect 21097 28917 21131 28951
rect 2789 28713 2823 28747
rect 11805 28713 11839 28747
rect 11989 28713 12023 28747
rect 16957 28713 16991 28747
rect 26617 28713 26651 28747
rect 28181 28713 28215 28747
rect 38209 28713 38243 28747
rect 20085 28645 20119 28679
rect 31217 28645 31251 28679
rect 4445 28577 4479 28611
rect 5641 28577 5675 28611
rect 8125 28577 8159 28611
rect 28273 28577 28307 28611
rect 30021 28577 30055 28611
rect 37657 28577 37691 28611
rect 1961 28509 1995 28543
rect 2881 28509 2915 28543
rect 4261 28509 4295 28543
rect 8217 28509 8251 28543
rect 15669 28509 15703 28543
rect 18521 28509 18555 28543
rect 20361 28509 20395 28543
rect 20821 28509 20855 28543
rect 20913 28509 20947 28543
rect 21097 28509 21131 28543
rect 21189 28509 21223 28543
rect 21833 28509 21867 28543
rect 25237 28509 25271 28543
rect 27997 28509 28031 28543
rect 29837 28509 29871 28543
rect 31677 28509 31711 28543
rect 35817 28509 35851 28543
rect 38117 28509 38151 28543
rect 12173 28441 12207 28475
rect 18705 28441 18739 28475
rect 20085 28441 20119 28475
rect 21373 28441 21407 28475
rect 22078 28441 22112 28475
rect 25504 28441 25538 28475
rect 31033 28441 31067 28475
rect 31769 28441 31803 28475
rect 36001 28441 36035 28475
rect 8585 28373 8619 28407
rect 11973 28373 12007 28407
rect 20269 28373 20303 28407
rect 23213 28373 23247 28407
rect 27813 28373 27847 28407
rect 12265 28169 12299 28203
rect 15209 28169 15243 28203
rect 23565 28169 23599 28203
rect 29285 28169 29319 28203
rect 32321 28169 32355 28203
rect 35265 28169 35299 28203
rect 36001 28169 36035 28203
rect 17017 28101 17051 28135
rect 17233 28101 17267 28135
rect 20545 28101 20579 28135
rect 23765 28101 23799 28135
rect 24593 28101 24627 28135
rect 30389 28101 30423 28135
rect 1869 28033 1903 28067
rect 4353 28033 4387 28067
rect 8861 28033 8895 28067
rect 11897 28033 11931 28067
rect 13277 28033 13311 28067
rect 14749 28033 14783 28067
rect 15209 28033 15243 28067
rect 15945 28033 15979 28067
rect 16037 28033 16071 28067
rect 16129 28033 16163 28067
rect 16313 28033 16347 28067
rect 19717 28033 19751 28067
rect 19993 28033 20027 28067
rect 22753 28033 22787 28067
rect 22937 28033 22971 28067
rect 24409 28033 24443 28067
rect 26157 28033 26191 28067
rect 28172 28033 28206 28067
rect 30113 28033 30147 28067
rect 30205 28033 30239 28067
rect 30941 28033 30975 28067
rect 31033 28033 31067 28067
rect 31217 28033 31251 28067
rect 32505 28033 32539 28067
rect 35081 28033 35115 28067
rect 35909 28033 35943 28067
rect 2053 27965 2087 27999
rect 2789 27965 2823 27999
rect 8769 27965 8803 27999
rect 11805 27965 11839 27999
rect 13369 27965 13403 27999
rect 15025 27965 15059 27999
rect 19901 27965 19935 27999
rect 21005 27965 21039 27999
rect 26249 27965 26283 27999
rect 27905 27965 27939 27999
rect 30389 27965 30423 27999
rect 31125 27965 31159 27999
rect 32689 27965 32723 27999
rect 12909 27897 12943 27931
rect 15669 27897 15703 27931
rect 19809 27897 19843 27931
rect 20821 27897 20855 27931
rect 9137 27829 9171 27863
rect 14887 27829 14921 27863
rect 16865 27829 16899 27863
rect 17049 27829 17083 27863
rect 19533 27829 19567 27863
rect 22845 27829 22879 27863
rect 23397 27829 23431 27863
rect 23581 27829 23615 27863
rect 24225 27829 24259 27863
rect 25789 27829 25823 27863
rect 31401 27829 31435 27863
rect 37565 27829 37599 27863
rect 2145 27625 2179 27659
rect 15945 27625 15979 27659
rect 19901 27625 19935 27659
rect 21005 27625 21039 27659
rect 30573 27625 30607 27659
rect 31769 27625 31803 27659
rect 9873 27557 9907 27591
rect 11161 27557 11195 27591
rect 13369 27557 13403 27591
rect 27537 27557 27571 27591
rect 28549 27557 28583 27591
rect 9597 27489 9631 27523
rect 10885 27489 10919 27523
rect 13093 27489 13127 27523
rect 18429 27489 18463 27523
rect 19441 27489 19475 27523
rect 23581 27489 23615 27523
rect 27445 27489 27479 27523
rect 31309 27489 31343 27523
rect 32321 27489 32355 27523
rect 36461 27489 36495 27523
rect 2237 27421 2271 27455
rect 9505 27421 9539 27455
rect 10793 27421 10827 27455
rect 13001 27421 13035 27455
rect 15393 27421 15427 27455
rect 15485 27421 15519 27455
rect 15669 27421 15703 27455
rect 15761 27421 15795 27455
rect 19625 27421 19659 27455
rect 19993 27421 20027 27455
rect 23029 27421 23063 27455
rect 23121 27421 23155 27455
rect 24041 27421 24075 27455
rect 25145 27421 25179 27455
rect 25329 27421 25363 27455
rect 27353 27421 27387 27455
rect 27629 27421 27663 27455
rect 28733 27421 28767 27455
rect 30573 27421 30607 27455
rect 30757 27421 30791 27455
rect 31401 27421 31435 27455
rect 32229 27421 32263 27455
rect 32413 27421 32447 27455
rect 18162 27353 18196 27387
rect 20821 27353 20855 27387
rect 22845 27353 22879 27387
rect 36645 27353 36679 27387
rect 38301 27353 38335 27387
rect 17049 27285 17083 27319
rect 21021 27285 21055 27319
rect 21189 27285 21223 27319
rect 22943 27285 22977 27319
rect 23857 27285 23891 27319
rect 23949 27285 23983 27319
rect 25329 27285 25363 27319
rect 27169 27285 27203 27319
rect 18245 27081 18279 27115
rect 19073 27081 19107 27115
rect 25697 27081 25731 27115
rect 37565 27081 37599 27115
rect 17417 27013 17451 27047
rect 4261 26945 4295 26979
rect 8585 26945 8619 26979
rect 8769 26945 8803 26979
rect 9229 26945 9263 26979
rect 9413 26945 9447 26979
rect 11713 26945 11747 26979
rect 11897 26945 11931 26979
rect 12449 26945 12483 26979
rect 12633 26945 12667 26979
rect 12817 26945 12851 26979
rect 18061 26945 18095 26979
rect 19073 26945 19107 26979
rect 23489 26945 23523 26979
rect 24317 26945 24351 26979
rect 24501 26945 24535 26979
rect 25513 26945 25547 26979
rect 25789 26945 25823 26979
rect 26249 26945 26283 26979
rect 26433 26945 26467 26979
rect 29837 26945 29871 26979
rect 37473 26945 37507 26979
rect 8677 26877 8711 26911
rect 19349 26877 19383 26911
rect 23581 26877 23615 26911
rect 29561 26877 29595 26911
rect 17049 26809 17083 26843
rect 17601 26809 17635 26843
rect 19165 26809 19199 26843
rect 25513 26809 25547 26843
rect 4077 26741 4111 26775
rect 9413 26741 9447 26775
rect 11805 26741 11839 26775
rect 17417 26741 17451 26775
rect 23489 26741 23523 26775
rect 23857 26741 23891 26775
rect 24409 26741 24443 26775
rect 26341 26741 26375 26775
rect 8585 26537 8619 26571
rect 9597 26537 9631 26571
rect 12817 26537 12851 26571
rect 17417 26537 17451 26571
rect 22569 26537 22603 26571
rect 25789 26537 25823 26571
rect 26157 26537 26191 26571
rect 26617 26537 26651 26571
rect 26801 26537 26835 26571
rect 27813 26537 27847 26571
rect 27997 26537 28031 26571
rect 11069 26469 11103 26503
rect 15577 26469 15611 26503
rect 19717 26469 19751 26503
rect 24869 26469 24903 26503
rect 29837 26469 29871 26503
rect 3985 26401 4019 26435
rect 4445 26401 4479 26435
rect 9413 26401 9447 26435
rect 14565 26401 14599 26435
rect 15945 26401 15979 26435
rect 16037 26401 16071 26435
rect 26065 26401 26099 26435
rect 8309 26333 8343 26367
rect 8401 26333 8435 26367
rect 9321 26333 9355 26367
rect 10793 26333 10827 26367
rect 10885 26333 10919 26367
rect 11989 26333 12023 26367
rect 12173 26333 12207 26367
rect 14289 26333 14323 26367
rect 15761 26333 15795 26367
rect 15853 26333 15887 26367
rect 17601 26333 17635 26367
rect 17877 26333 17911 26367
rect 19441 26333 19475 26367
rect 21189 26333 21223 26367
rect 23765 26333 23799 26367
rect 24041 26333 24075 26367
rect 24593 26333 24627 26367
rect 24685 26333 24719 26367
rect 26157 26333 26191 26367
rect 27721 26333 27755 26367
rect 27905 26333 27939 26367
rect 28181 26333 28215 26367
rect 29009 26333 29043 26367
rect 29193 26333 29227 26367
rect 30021 26333 30055 26367
rect 4169 26265 4203 26299
rect 11069 26265 11103 26299
rect 12081 26265 12115 26299
rect 12785 26265 12819 26299
rect 13001 26265 13035 26299
rect 19717 26265 19751 26299
rect 21456 26265 21490 26299
rect 24869 26265 24903 26299
rect 26985 26265 27019 26299
rect 12633 26197 12667 26231
rect 17785 26197 17819 26231
rect 19533 26197 19567 26231
rect 26775 26197 26809 26231
rect 27445 26197 27479 26231
rect 29101 26197 29135 26231
rect 8585 25993 8619 26027
rect 11805 25993 11839 26027
rect 13829 25993 13863 26027
rect 15853 25993 15887 26027
rect 17233 25993 17267 26027
rect 17401 25993 17435 26027
rect 25697 25993 25731 26027
rect 8769 25925 8803 25959
rect 8953 25925 8987 25959
rect 9505 25925 9539 25959
rect 17601 25925 17635 25959
rect 18153 25925 18187 25959
rect 20646 25925 20680 25959
rect 25881 25925 25915 25959
rect 29000 25925 29034 25959
rect 9413 25857 9447 25891
rect 9597 25857 9631 25891
rect 11713 25857 11747 25891
rect 11897 25857 11931 25891
rect 12449 25857 12483 25891
rect 12716 25857 12750 25891
rect 15761 25857 15795 25891
rect 20913 25857 20947 25891
rect 23397 25857 23431 25891
rect 25605 25857 25639 25891
rect 26433 25857 26467 25891
rect 27445 25857 27479 25891
rect 27537 25857 27571 25891
rect 27721 25857 27755 25891
rect 27813 25857 27847 25891
rect 30757 25857 30791 25891
rect 37473 25857 37507 25891
rect 14841 25789 14875 25823
rect 15301 25789 15335 25823
rect 28733 25789 28767 25823
rect 30665 25789 30699 25823
rect 15117 25721 15151 25755
rect 18337 25721 18371 25755
rect 24685 25721 24719 25755
rect 30113 25721 30147 25755
rect 17417 25653 17451 25687
rect 19533 25653 19567 25687
rect 25881 25653 25915 25687
rect 26525 25653 26559 25687
rect 27261 25653 27295 25687
rect 31125 25653 31159 25687
rect 37565 25653 37599 25687
rect 38301 25653 38335 25687
rect 4077 25449 4111 25483
rect 12725 25449 12759 25483
rect 14933 25449 14967 25483
rect 15301 25449 15335 25483
rect 18061 25449 18095 25483
rect 19717 25449 19751 25483
rect 23765 25449 23799 25483
rect 24593 25449 24627 25483
rect 27537 25381 27571 25415
rect 19625 25313 19659 25347
rect 22385 25313 22419 25347
rect 27353 25313 27387 25347
rect 30849 25313 30883 25347
rect 37841 25313 37875 25347
rect 38117 25313 38151 25347
rect 38301 25313 38335 25347
rect 3985 25245 4019 25279
rect 12909 25245 12943 25279
rect 14841 25245 14875 25279
rect 18061 25245 18095 25279
rect 18245 25245 18279 25279
rect 19809 25245 19843 25279
rect 19901 25245 19935 25279
rect 21465 25245 21499 25279
rect 24777 25245 24811 25279
rect 24869 25245 24903 25279
rect 27077 25245 27111 25279
rect 27169 25245 27203 25279
rect 27261 25245 27295 25279
rect 30573 25245 30607 25279
rect 30665 25245 30699 25279
rect 31309 25245 31343 25279
rect 31493 25245 31527 25279
rect 17233 25177 17267 25211
rect 17417 25177 17451 25211
rect 22630 25177 22664 25211
rect 24593 25177 24627 25211
rect 17601 25109 17635 25143
rect 21281 25109 21315 25143
rect 30573 25109 30607 25143
rect 31401 25109 31435 25143
rect 26341 24905 26375 24939
rect 30021 24905 30055 24939
rect 31309 24905 31343 24939
rect 9413 24837 9447 24871
rect 24685 24837 24719 24871
rect 24885 24837 24919 24871
rect 25881 24837 25915 24871
rect 9643 24803 9677 24837
rect 25651 24803 25685 24837
rect 10241 24769 10275 24803
rect 16037 24769 16071 24803
rect 17601 24769 17635 24803
rect 17785 24769 17819 24803
rect 18245 24769 18279 24803
rect 18429 24769 18463 24803
rect 19901 24769 19935 24803
rect 20085 24769 20119 24803
rect 20729 24769 20763 24803
rect 21189 24769 21223 24803
rect 22845 24769 22879 24803
rect 26617 24769 26651 24803
rect 27353 24769 27387 24803
rect 27537 24769 27571 24803
rect 28089 24769 28123 24803
rect 28273 24769 28307 24803
rect 29101 24769 29135 24803
rect 29285 24769 29319 24803
rect 29962 24769 29996 24803
rect 30481 24769 30515 24803
rect 31125 24769 31159 24803
rect 31401 24769 31435 24803
rect 37473 24769 37507 24803
rect 3893 24701 3927 24735
rect 4077 24701 4111 24735
rect 5457 24701 5491 24735
rect 14197 24701 14231 24735
rect 14381 24701 14415 24735
rect 20637 24701 20671 24735
rect 22569 24701 22603 24735
rect 26341 24701 26375 24735
rect 27629 24701 27663 24735
rect 28181 24701 28215 24735
rect 9781 24633 9815 24667
rect 17417 24633 17451 24667
rect 20085 24633 20119 24667
rect 29837 24633 29871 24667
rect 9597 24565 9631 24599
rect 10425 24565 10459 24599
rect 18245 24565 18279 24599
rect 21373 24565 21407 24599
rect 24869 24565 24903 24599
rect 25053 24565 25087 24599
rect 25513 24565 25547 24599
rect 25697 24565 25731 24599
rect 26525 24565 26559 24599
rect 27169 24565 27203 24599
rect 29193 24565 29227 24599
rect 30389 24565 30423 24599
rect 30941 24565 30975 24599
rect 37565 24565 37599 24599
rect 38301 24565 38335 24599
rect 4077 24361 4111 24395
rect 9229 24361 9263 24395
rect 11713 24361 11747 24395
rect 13737 24361 13771 24395
rect 22477 24361 22511 24395
rect 25053 24361 25087 24395
rect 26525 24361 26559 24395
rect 26709 24361 26743 24395
rect 28917 24361 28951 24395
rect 29745 24361 29779 24395
rect 23673 24293 23707 24327
rect 18705 24225 18739 24259
rect 25145 24225 25179 24259
rect 26801 24225 26835 24259
rect 27813 24225 27847 24259
rect 28457 24225 28491 24259
rect 28641 24225 28675 24259
rect 37841 24225 37875 24259
rect 38117 24225 38151 24259
rect 38301 24225 38335 24259
rect 3985 24157 4019 24191
rect 8585 24157 8619 24191
rect 9413 24157 9447 24191
rect 10333 24157 10367 24191
rect 13001 24157 13035 24191
rect 13553 24157 13587 24191
rect 14749 24157 14783 24191
rect 16966 24157 17000 24191
rect 17509 24157 17543 24191
rect 17693 24157 17727 24191
rect 17785 24157 17819 24191
rect 17923 24157 17957 24191
rect 18613 24157 18647 24191
rect 18797 24157 18831 24191
rect 22753 24157 22787 24191
rect 22842 24154 22876 24188
rect 22942 24157 22976 24191
rect 23121 24157 23155 24191
rect 23581 24157 23615 24191
rect 23765 24157 23799 24191
rect 24869 24157 24903 24191
rect 26893 24157 26927 24191
rect 27721 24157 27755 24191
rect 27905 24157 27939 24191
rect 28549 24157 28583 24191
rect 28733 24157 28767 24191
rect 29929 24157 29963 24191
rect 30205 24157 30239 24191
rect 9597 24089 9631 24123
rect 10578 24089 10612 24123
rect 15016 24089 15050 24123
rect 16681 24089 16715 24123
rect 20269 24089 20303 24123
rect 8493 24021 8527 24055
rect 12909 24021 12943 24055
rect 16129 24021 16163 24055
rect 16779 24021 16813 24055
rect 16865 24021 16899 24055
rect 18153 24021 18187 24055
rect 21557 24021 21591 24055
rect 24685 24021 24719 24055
rect 30113 24021 30147 24055
rect 14105 23817 14139 23851
rect 20453 23817 20487 23851
rect 22201 23817 22235 23851
rect 29193 23817 29227 23851
rect 10041 23749 10075 23783
rect 10241 23749 10275 23783
rect 12265 23749 12299 23783
rect 17325 23749 17359 23783
rect 19450 23749 19484 23783
rect 20913 23749 20947 23783
rect 23581 23749 23615 23783
rect 23765 23749 23799 23783
rect 29377 23749 29411 23783
rect 29561 23749 29595 23783
rect 35725 23749 35759 23783
rect 9045 23681 9079 23715
rect 9229 23681 9263 23715
rect 9413 23681 9447 23715
rect 13277 23681 13311 23715
rect 13369 23681 13403 23715
rect 14289 23681 14323 23715
rect 14749 23681 14783 23715
rect 17233 23681 17267 23715
rect 17509 23681 17543 23715
rect 22109 23681 22143 23715
rect 22845 23681 22879 23715
rect 24768 23681 24802 23715
rect 28365 23681 28399 23715
rect 33885 23681 33919 23715
rect 12449 23613 12483 23647
rect 14381 23613 14415 23647
rect 19717 23613 19751 23647
rect 24501 23613 24535 23647
rect 28273 23613 28307 23647
rect 28733 23613 28767 23647
rect 34069 23613 34103 23647
rect 9045 23545 9079 23579
rect 13645 23545 13679 23579
rect 17509 23545 17543 23579
rect 20637 23545 20671 23579
rect 9137 23477 9171 23511
rect 9873 23477 9907 23511
rect 10057 23477 10091 23511
rect 13461 23477 13495 23511
rect 14289 23477 14323 23511
rect 18337 23477 18371 23511
rect 22937 23477 22971 23511
rect 25881 23477 25915 23511
rect 10149 23273 10183 23307
rect 14381 23273 14415 23307
rect 17049 23273 17083 23307
rect 20361 23273 20395 23307
rect 33885 23273 33919 23307
rect 17233 23205 17267 23239
rect 20177 23205 20211 23239
rect 26801 23205 26835 23239
rect 31033 23205 31067 23239
rect 18153 23137 18187 23171
rect 20453 23137 20487 23171
rect 26341 23137 26375 23171
rect 30573 23137 30607 23171
rect 31769 23137 31803 23171
rect 2329 23069 2363 23103
rect 2973 23069 3007 23103
rect 9413 23069 9447 23103
rect 9597 23069 9631 23103
rect 10057 23069 10091 23103
rect 10241 23069 10275 23103
rect 10793 23069 10827 23103
rect 11049 23069 11083 23103
rect 12725 23069 12759 23103
rect 12909 23069 12943 23103
rect 14289 23069 14323 23103
rect 16221 23069 16255 23103
rect 17785 23069 17819 23103
rect 17969 23069 18003 23103
rect 20545 23069 20579 23103
rect 21465 23069 21499 23103
rect 21925 23069 21959 23103
rect 22937 23069 22971 23103
rect 23489 23069 23523 23103
rect 23673 23069 23707 23103
rect 26433 23069 26467 23103
rect 30665 23069 30699 23103
rect 31861 23069 31895 23103
rect 33793 23069 33827 23103
rect 37841 23069 37875 23103
rect 16405 23001 16439 23035
rect 16865 23001 16899 23035
rect 18705 23001 18739 23035
rect 22109 23001 22143 23035
rect 22293 23001 22327 23035
rect 2237 22933 2271 22967
rect 9505 22933 9539 22967
rect 12173 22933 12207 22967
rect 12909 22933 12943 22967
rect 17065 22933 17099 22967
rect 18797 22933 18831 22967
rect 21281 22933 21315 22967
rect 22753 22933 22787 22967
rect 23673 22933 23707 22967
rect 31493 22933 31527 22967
rect 12633 22729 12667 22763
rect 15485 22729 15519 22763
rect 17233 22729 17267 22763
rect 18245 22729 18279 22763
rect 18429 22729 18463 22763
rect 30573 22729 30607 22763
rect 3525 22661 3559 22695
rect 15117 22661 15151 22695
rect 22468 22661 22502 22695
rect 24777 22661 24811 22695
rect 3709 22593 3743 22627
rect 8953 22593 8987 22627
rect 12817 22593 12851 22627
rect 15301 22593 15335 22627
rect 15933 22593 15967 22627
rect 16037 22593 16071 22627
rect 16865 22593 16899 22627
rect 17049 22593 17083 22627
rect 18370 22593 18404 22627
rect 20453 22593 20487 22627
rect 20545 22593 20579 22627
rect 20729 22593 20763 22627
rect 22201 22593 22235 22627
rect 30514 22593 30548 22627
rect 31033 22593 31067 22627
rect 37473 22593 37507 22627
rect 1869 22525 1903 22559
rect 9045 22525 9079 22559
rect 9321 22525 9355 22559
rect 18889 22525 18923 22559
rect 30941 22525 30975 22559
rect 23581 22457 23615 22491
rect 24961 22457 24995 22491
rect 15945 22389 15979 22423
rect 16313 22389 16347 22423
rect 16865 22389 16899 22423
rect 18797 22389 18831 22423
rect 20913 22389 20947 22423
rect 30389 22389 30423 22423
rect 37565 22389 37599 22423
rect 13369 22185 13403 22219
rect 13737 22185 13771 22219
rect 14933 22185 14967 22219
rect 15577 22185 15611 22219
rect 20177 22185 20211 22219
rect 20821 22185 20855 22219
rect 31125 22185 31159 22219
rect 2789 22049 2823 22083
rect 12817 22049 12851 22083
rect 14749 22049 14783 22083
rect 15669 22049 15703 22083
rect 17417 22049 17451 22083
rect 17877 22049 17911 22083
rect 27353 22049 27387 22083
rect 37197 22049 37231 22083
rect 38117 22049 38151 22083
rect 38301 22049 38335 22083
rect 1593 21981 1627 22015
rect 10701 21981 10735 22015
rect 13369 21981 13403 22015
rect 13461 21981 13495 22015
rect 14933 21981 14967 22015
rect 15853 21981 15887 22015
rect 17325 21981 17359 22015
rect 20085 21981 20119 22015
rect 20269 21981 20303 22015
rect 21097 21981 21131 22015
rect 23673 21981 23707 22015
rect 23857 21981 23891 22015
rect 24869 21981 24903 22015
rect 26893 21981 26927 22015
rect 27077 21981 27111 22015
rect 27169 21981 27203 22015
rect 27445 21981 27479 22015
rect 29745 21981 29779 22015
rect 1777 21913 1811 21947
rect 10946 21913 10980 21947
rect 12633 21913 12667 21947
rect 14473 21913 14507 21947
rect 15577 21913 15611 21947
rect 25114 21913 25148 21947
rect 29990 21913 30024 21947
rect 12081 21845 12115 21879
rect 15117 21845 15151 21879
rect 16037 21845 16071 21879
rect 17693 21845 17727 21879
rect 23857 21845 23891 21879
rect 26249 21845 26283 21879
rect 2421 21641 2455 21675
rect 14013 21641 14047 21675
rect 15117 21641 15151 21675
rect 21005 21641 21039 21675
rect 21373 21641 21407 21675
rect 24409 21641 24443 21675
rect 29653 21641 29687 21675
rect 9045 21573 9079 21607
rect 12081 21573 12115 21607
rect 12725 21573 12759 21607
rect 17325 21573 17359 21607
rect 17509 21573 17543 21607
rect 35449 21573 35483 21607
rect 1685 21505 1719 21539
rect 2513 21505 2547 21539
rect 2973 21505 3007 21539
rect 8769 21505 8803 21539
rect 8861 21505 8895 21539
rect 9505 21505 9539 21539
rect 9689 21505 9723 21539
rect 11897 21505 11931 21539
rect 13185 21505 13219 21539
rect 13921 21505 13955 21539
rect 14105 21505 14139 21539
rect 14565 21505 14599 21539
rect 15577 21505 15611 21539
rect 15853 21505 15887 21539
rect 18797 21505 18831 21539
rect 18981 21505 19015 21539
rect 20913 21505 20947 21539
rect 21189 21505 21223 21539
rect 22661 21505 22695 21539
rect 23765 21505 23799 21539
rect 23949 21505 23983 21539
rect 24041 21505 24075 21539
rect 24133 21505 24167 21539
rect 27721 21505 27755 21539
rect 27988 21505 28022 21539
rect 29561 21505 29595 21539
rect 29745 21505 29779 21539
rect 32965 21505 32999 21539
rect 33609 21505 33643 21539
rect 9045 21437 9079 21471
rect 13001 21437 13035 21471
rect 14841 21437 14875 21471
rect 15669 21437 15703 21471
rect 22753 21437 22787 21471
rect 33057 21437 33091 21471
rect 33793 21437 33827 21471
rect 15577 21369 15611 21403
rect 17693 21369 17727 21403
rect 23029 21369 23063 21403
rect 3065 21301 3099 21335
rect 9689 21301 9723 21335
rect 12265 21301 12299 21335
rect 13185 21301 13219 21335
rect 13369 21301 13403 21335
rect 14933 21301 14967 21335
rect 17509 21301 17543 21335
rect 18889 21301 18923 21335
rect 29101 21301 29135 21335
rect 8401 21097 8435 21131
rect 9137 21097 9171 21131
rect 13553 21097 13587 21131
rect 17141 21097 17175 21131
rect 27997 21097 28031 21131
rect 14841 21029 14875 21063
rect 1593 20961 1627 20995
rect 3249 20961 3283 20995
rect 8585 20961 8619 20995
rect 9505 20961 9539 20995
rect 14565 20961 14599 20995
rect 14657 20961 14691 20995
rect 22569 20961 22603 20995
rect 24593 20961 24627 20995
rect 26433 20961 26467 20995
rect 26709 20961 26743 20995
rect 3433 20893 3467 20927
rect 8309 20893 8343 20927
rect 9321 20893 9355 20927
rect 10333 20893 10367 20927
rect 12173 20893 12207 20927
rect 14381 20893 14415 20927
rect 14473 20893 14507 20927
rect 17233 20893 17267 20927
rect 17877 20893 17911 20927
rect 18061 20893 18095 20927
rect 18521 20893 18555 20927
rect 19625 20893 19659 20927
rect 20821 20893 20855 20927
rect 24849 20893 24883 20927
rect 27721 20893 27755 20927
rect 28457 20893 28491 20927
rect 28641 20893 28675 20927
rect 10578 20825 10612 20859
rect 12440 20825 12474 20859
rect 18705 20825 18739 20859
rect 19809 20825 19843 20859
rect 27997 20825 28031 20859
rect 8585 20757 8619 20791
rect 11713 20757 11747 20791
rect 17969 20757 18003 20791
rect 18889 20757 18923 20791
rect 19441 20757 19475 20791
rect 25973 20757 26007 20791
rect 27813 20757 27847 20791
rect 28457 20757 28491 20791
rect 8969 20553 9003 20587
rect 9689 20553 9723 20587
rect 13645 20553 13679 20587
rect 16957 20553 16991 20587
rect 20085 20553 20119 20587
rect 27337 20553 27371 20587
rect 30573 20553 30607 20587
rect 1961 20485 1995 20519
rect 8769 20485 8803 20519
rect 19165 20485 19199 20519
rect 19257 20485 19291 20519
rect 27537 20485 27571 20519
rect 27997 20485 28031 20519
rect 9597 20417 9631 20451
rect 9781 20417 9815 20451
rect 12817 20417 12851 20451
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 14933 20417 14967 20451
rect 16865 20417 16899 20451
rect 17693 20417 17727 20451
rect 18981 20417 19015 20451
rect 19349 20417 19383 20451
rect 21198 20417 21232 20451
rect 21465 20417 21499 20451
rect 22293 20417 22327 20451
rect 26341 20417 26375 20451
rect 26433 20417 26467 20451
rect 26617 20417 26651 20451
rect 28181 20417 28215 20451
rect 28273 20417 28307 20451
rect 30514 20417 30548 20451
rect 31493 20417 31527 20451
rect 3617 20349 3651 20383
rect 3801 20349 3835 20383
rect 22385 20349 22419 20383
rect 25973 20349 26007 20383
rect 31033 20349 31067 20383
rect 9137 20281 9171 20315
rect 12633 20281 12667 20315
rect 19533 20281 19567 20315
rect 22661 20281 22695 20315
rect 31585 20281 31619 20315
rect 8953 20213 8987 20247
rect 13461 20213 13495 20247
rect 15025 20213 15059 20247
rect 17601 20213 17635 20247
rect 27169 20213 27203 20247
rect 27353 20213 27387 20247
rect 27997 20213 28031 20247
rect 30389 20213 30423 20247
rect 30941 20213 30975 20247
rect 2697 20009 2731 20043
rect 3433 20009 3467 20043
rect 18337 20009 18371 20043
rect 20637 20009 20671 20043
rect 21281 20009 21315 20043
rect 26433 20009 26467 20043
rect 27169 20009 27203 20043
rect 31125 20009 31159 20043
rect 31677 20009 31711 20043
rect 2145 19941 2179 19975
rect 27353 19941 27387 19975
rect 27905 19941 27939 19975
rect 15301 19873 15335 19907
rect 17135 19873 17169 19907
rect 17233 19873 17267 19907
rect 30665 19873 30699 19907
rect 31861 19873 31895 19907
rect 2789 19805 2823 19839
rect 14289 19805 14323 19839
rect 15209 19805 15243 19839
rect 16853 19795 16887 19829
rect 17049 19805 17083 19839
rect 17417 19805 17451 19839
rect 18705 19805 18739 19839
rect 20269 19805 20303 19839
rect 21465 19805 21499 19839
rect 23673 19805 23707 19839
rect 24041 19805 24075 19839
rect 26065 19805 26099 19839
rect 26249 19805 26283 19839
rect 26985 19805 27019 19839
rect 27169 19805 27203 19839
rect 27813 19805 27847 19839
rect 27997 19805 28031 19839
rect 29745 19805 29779 19839
rect 29929 19805 29963 19839
rect 30757 19805 30791 19839
rect 31953 19805 31987 19839
rect 37473 19805 37507 19839
rect 16129 19737 16163 19771
rect 18889 19737 18923 19771
rect 23765 19737 23799 19771
rect 23857 19737 23891 19771
rect 14473 19669 14507 19703
rect 15577 19669 15611 19703
rect 16221 19669 16255 19703
rect 17601 19669 17635 19703
rect 18521 19669 18555 19703
rect 18613 19669 18647 19703
rect 20637 19669 20671 19703
rect 20821 19669 20855 19703
rect 23489 19669 23523 19703
rect 29837 19669 29871 19703
rect 37565 19669 37599 19703
rect 13553 19465 13587 19499
rect 17141 19465 17175 19499
rect 18337 19465 18371 19499
rect 20085 19465 20119 19499
rect 30113 19465 30147 19499
rect 2789 19397 2823 19431
rect 10517 19397 10551 19431
rect 17693 19397 17727 19431
rect 19717 19397 19751 19431
rect 19933 19397 19967 19431
rect 27261 19397 27295 19431
rect 29000 19397 29034 19431
rect 2513 19329 2547 19363
rect 4077 19329 4111 19363
rect 9873 19329 9907 19363
rect 10057 19329 10091 19363
rect 10149 19329 10183 19363
rect 10241 19329 10275 19363
rect 12173 19329 12207 19363
rect 12429 19329 12463 19363
rect 14749 19329 14783 19363
rect 18429 19329 18463 19363
rect 20729 19329 20763 19363
rect 21005 19329 21039 19363
rect 22293 19329 22327 19363
rect 22477 19329 22511 19363
rect 22937 19329 22971 19363
rect 23949 19329 23983 19363
rect 24133 19329 24167 19363
rect 24225 19329 24259 19363
rect 24501 19329 24535 19363
rect 25789 19329 25823 19363
rect 25973 19329 26007 19363
rect 30573 19329 30607 19363
rect 3801 19261 3835 19295
rect 16957 19261 16991 19295
rect 17233 19261 17267 19295
rect 20821 19261 20855 19295
rect 20913 19261 20947 19295
rect 23213 19261 23247 19295
rect 24409 19261 24443 19295
rect 26157 19261 26191 19295
rect 28733 19261 28767 19295
rect 30849 19261 30883 19295
rect 14933 19193 14967 19227
rect 17693 19193 17727 19227
rect 20545 19193 20579 19227
rect 27445 19193 27479 19227
rect 19901 19125 19935 19159
rect 22385 19125 22419 19159
rect 23029 19125 23063 19159
rect 23489 19125 23523 19159
rect 37841 19125 37875 19159
rect 9413 18921 9447 18955
rect 10149 18921 10183 18955
rect 10333 18921 10367 18955
rect 12173 18921 12207 18955
rect 17785 18921 17819 18955
rect 20177 18921 20211 18955
rect 23489 18921 23523 18955
rect 31677 18921 31711 18955
rect 13553 18853 13587 18887
rect 22937 18853 22971 18887
rect 27445 18853 27479 18887
rect 31033 18853 31067 18887
rect 4813 18785 4847 18819
rect 17325 18785 17359 18819
rect 20545 18785 20579 18819
rect 25053 18785 25087 18819
rect 28273 18785 28307 18819
rect 31217 18785 31251 18819
rect 37841 18785 37875 18819
rect 38117 18785 38151 18819
rect 38301 18785 38335 18819
rect 2237 18717 2271 18751
rect 2789 18717 2823 18751
rect 9137 18717 9171 18751
rect 9229 18717 9263 18751
rect 9505 18717 9539 18751
rect 10793 18717 10827 18751
rect 11060 18717 11094 18751
rect 13737 18717 13771 18751
rect 14289 18717 14323 18751
rect 16129 18717 16163 18751
rect 17049 18717 17083 18751
rect 17233 18717 17267 18751
rect 17417 18717 17451 18751
rect 17612 18717 17646 18751
rect 20453 18717 20487 18751
rect 20637 18717 20671 18751
rect 20913 18717 20947 18751
rect 22201 18717 22235 18751
rect 23121 18717 23155 18751
rect 24961 18717 24995 18751
rect 27629 18717 27663 18751
rect 28457 18717 28491 18751
rect 28549 18717 28583 18751
rect 31677 18717 31711 18751
rect 31861 18717 31895 18751
rect 2053 18649 2087 18683
rect 3341 18649 3375 18683
rect 3985 18649 4019 18683
rect 9965 18649 9999 18683
rect 14556 18649 14590 18683
rect 22385 18649 22419 18683
rect 30757 18649 30791 18683
rect 9321 18581 9355 18615
rect 10165 18581 10199 18615
rect 15669 18581 15703 18615
rect 16221 18581 16255 18615
rect 20821 18581 20855 18615
rect 23213 18581 23247 18615
rect 23305 18581 23339 18615
rect 24593 18581 24627 18615
rect 28273 18581 28307 18615
rect 10425 18377 10459 18411
rect 12357 18377 12391 18411
rect 16865 18377 16899 18411
rect 20637 18377 20671 18411
rect 22569 18377 22603 18411
rect 23213 18377 23247 18411
rect 31677 18377 31711 18411
rect 4445 18309 4479 18343
rect 9873 18309 9907 18343
rect 13001 18309 13035 18343
rect 14749 18309 14783 18343
rect 17233 18309 17267 18343
rect 18705 18309 18739 18343
rect 25789 18309 25823 18343
rect 25973 18309 26007 18343
rect 4169 18241 4203 18275
rect 8861 18241 8895 18275
rect 8953 18241 8987 18275
rect 9597 18241 9631 18275
rect 10333 18241 10367 18275
rect 10517 18241 10551 18275
rect 12265 18241 12299 18275
rect 12541 18241 12575 18275
rect 15761 18241 15795 18275
rect 16037 18241 16071 18275
rect 16129 18241 16163 18275
rect 16313 18241 16347 18275
rect 17003 18241 17037 18275
rect 17141 18241 17175 18275
rect 17361 18241 17395 18275
rect 17509 18241 17543 18275
rect 20361 18241 20395 18275
rect 22201 18241 22235 18275
rect 23397 18241 23431 18275
rect 23489 18241 23523 18275
rect 23673 18241 23707 18275
rect 27261 18241 27295 18275
rect 27445 18241 27479 18275
rect 27537 18241 27571 18275
rect 27997 18241 28031 18275
rect 28253 18241 28287 18275
rect 30481 18241 30515 18275
rect 30665 18241 30699 18275
rect 30941 18241 30975 18275
rect 31585 18241 31619 18275
rect 31769 18241 31803 18275
rect 32321 18241 32355 18275
rect 32505 18241 32539 18275
rect 1869 18173 1903 18207
rect 2053 18173 2087 18207
rect 2789 18173 2823 18207
rect 9873 18173 9907 18207
rect 20637 18173 20671 18207
rect 22293 18173 22327 18207
rect 15853 18105 15887 18139
rect 27261 18105 27295 18139
rect 9137 18037 9171 18071
rect 9689 18037 9723 18071
rect 12541 18037 12575 18071
rect 18797 18037 18831 18071
rect 20453 18037 20487 18071
rect 23581 18037 23615 18071
rect 26157 18037 26191 18071
rect 29377 18037 29411 18071
rect 31125 18037 31159 18071
rect 32321 18037 32355 18071
rect 37473 18037 37507 18071
rect 1777 17833 1811 17867
rect 2329 17833 2363 17867
rect 9229 17833 9263 17867
rect 13093 17833 13127 17867
rect 14565 17833 14599 17867
rect 18153 17833 18187 17867
rect 27537 17833 27571 17867
rect 28089 17833 28123 17867
rect 32045 17833 32079 17867
rect 9321 17765 9355 17799
rect 20361 17765 20395 17799
rect 31861 17765 31895 17799
rect 9413 17697 9447 17731
rect 18613 17697 18647 17731
rect 20085 17697 20119 17731
rect 30849 17697 30883 17731
rect 31033 17697 31067 17731
rect 36461 17697 36495 17731
rect 38301 17697 38335 17731
rect 2421 17629 2455 17663
rect 3065 17629 3099 17663
rect 3985 17629 4019 17663
rect 4261 17629 4295 17663
rect 9137 17629 9171 17663
rect 9873 17629 9907 17663
rect 10057 17629 10091 17663
rect 11713 17629 11747 17663
rect 14841 17629 14875 17663
rect 14933 17629 14967 17663
rect 15025 17629 15059 17663
rect 15209 17629 15243 17663
rect 18521 17629 18555 17663
rect 19993 17629 20027 17663
rect 25973 17629 26007 17663
rect 26341 17629 26375 17663
rect 26433 17629 26467 17663
rect 27445 17629 27479 17663
rect 27629 17629 27663 17663
rect 28273 17629 28307 17663
rect 28549 17629 28583 17663
rect 30757 17629 30791 17663
rect 30941 17629 30975 17663
rect 9965 17561 9999 17595
rect 11958 17561 11992 17595
rect 15669 17561 15703 17595
rect 17417 17561 17451 17595
rect 22569 17561 22603 17595
rect 26065 17561 26099 17595
rect 26157 17561 26191 17595
rect 31585 17561 31619 17595
rect 36645 17561 36679 17595
rect 2973 17493 3007 17527
rect 21281 17493 21315 17527
rect 25789 17493 25823 17527
rect 28457 17493 28491 17527
rect 30573 17493 30607 17527
rect 23949 17289 23983 17323
rect 25957 17289 25991 17323
rect 27261 17289 27295 17323
rect 30297 17289 30331 17323
rect 37565 17289 37599 17323
rect 3525 17221 3559 17255
rect 17325 17221 17359 17255
rect 17693 17221 17727 17255
rect 21097 17221 21131 17255
rect 23121 17221 23155 17255
rect 26157 17221 26191 17255
rect 13001 17153 13035 17187
rect 13277 17153 13311 17187
rect 13829 17153 13863 17187
rect 14096 17153 14130 17187
rect 16062 17153 16096 17187
rect 17509 17153 17543 17187
rect 19441 17153 19475 17187
rect 21005 17153 21039 17187
rect 21189 17153 21223 17187
rect 22937 17153 22971 17187
rect 23213 17153 23247 17187
rect 23305 17153 23339 17187
rect 24317 17153 24351 17187
rect 25145 17153 25179 17187
rect 27169 17153 27203 17187
rect 27445 17153 27479 17187
rect 30113 17153 30147 17187
rect 30389 17153 30423 17187
rect 36921 17153 36955 17187
rect 37657 17153 37691 17187
rect 1869 17085 1903 17119
rect 3709 17085 3743 17119
rect 19533 17085 19567 17119
rect 24409 17085 24443 17119
rect 25329 17085 25363 17119
rect 27537 17085 27571 17119
rect 13093 17017 13127 17051
rect 13185 17017 13219 17051
rect 15209 17017 15243 17051
rect 19809 17017 19843 17051
rect 24961 17017 24995 17051
rect 25789 17017 25823 17051
rect 12817 16949 12851 16983
rect 16221 16949 16255 16983
rect 23489 16949 23523 16983
rect 25973 16949 26007 16983
rect 27353 16949 27387 16983
rect 30113 16949 30147 16983
rect 36829 16949 36863 16983
rect 38117 16949 38151 16983
rect 2145 16745 2179 16779
rect 12909 16745 12943 16779
rect 13461 16745 13495 16779
rect 14749 16745 14783 16779
rect 16865 16745 16899 16779
rect 17693 16745 17727 16779
rect 21005 16745 21039 16779
rect 21649 16745 21683 16779
rect 31217 16745 31251 16779
rect 10793 16677 10827 16711
rect 30297 16677 30331 16711
rect 9229 16609 9263 16643
rect 10517 16609 10551 16643
rect 11253 16609 11287 16643
rect 11805 16609 11839 16643
rect 14289 16609 14323 16643
rect 25789 16609 25823 16643
rect 26065 16609 26099 16643
rect 28365 16609 28399 16643
rect 36461 16609 36495 16643
rect 36645 16609 36679 16643
rect 38301 16609 38335 16643
rect 3433 16541 3467 16575
rect 4445 16541 4479 16575
rect 9321 16541 9355 16575
rect 10425 16541 10459 16575
rect 11529 16541 11563 16575
rect 12265 16541 12299 16575
rect 12403 16541 12437 16575
rect 12730 16541 12764 16575
rect 13369 16541 13403 16575
rect 13553 16541 13587 16575
rect 14381 16541 14415 16575
rect 14565 16541 14599 16575
rect 15853 16541 15887 16575
rect 16037 16541 16071 16575
rect 16957 16541 16991 16575
rect 17601 16541 17635 16575
rect 18245 16541 18279 16575
rect 18429 16541 18463 16575
rect 20637 16541 20671 16575
rect 21833 16541 21867 16575
rect 22109 16541 22143 16575
rect 28273 16541 28307 16575
rect 30665 16541 30699 16575
rect 31309 16541 31343 16575
rect 3157 16473 3191 16507
rect 4169 16473 4203 16507
rect 11621 16473 11655 16507
rect 12541 16473 12575 16507
rect 12633 16473 12667 16507
rect 9689 16405 9723 16439
rect 11437 16405 11471 16439
rect 15669 16405 15703 16439
rect 18245 16405 18279 16439
rect 21005 16405 21039 16439
rect 21189 16405 21223 16439
rect 22017 16405 22051 16439
rect 27905 16405 27939 16439
rect 30205 16405 30239 16439
rect 16865 16201 16899 16235
rect 23397 16201 23431 16235
rect 3157 16133 3191 16167
rect 4537 16133 4571 16167
rect 17141 16133 17175 16167
rect 2237 16065 2271 16099
rect 2421 16065 2455 16099
rect 2881 16065 2915 16099
rect 3801 16065 3835 16099
rect 5273 16065 5307 16099
rect 10425 16065 10459 16099
rect 15669 16065 15703 16099
rect 17049 16065 17083 16099
rect 17233 16065 17267 16099
rect 17417 16065 17451 16099
rect 18133 16065 18167 16099
rect 21281 16065 21315 16099
rect 22017 16065 22051 16099
rect 22273 16065 22307 16099
rect 25145 16065 25179 16099
rect 27629 16065 27663 16099
rect 27813 16065 27847 16099
rect 28089 16065 28123 16099
rect 28273 16065 28307 16099
rect 29193 16065 29227 16099
rect 31125 16065 31159 16099
rect 31309 16065 31343 16099
rect 36921 16065 36955 16099
rect 5825 15997 5859 16031
rect 10517 15997 10551 16031
rect 10793 15997 10827 16031
rect 17877 15997 17911 16031
rect 24869 15997 24903 16031
rect 28917 15997 28951 16031
rect 29009 15997 29043 16031
rect 29101 15997 29135 16031
rect 30205 15997 30239 16031
rect 30665 15997 30699 16031
rect 21465 15929 21499 15963
rect 30573 15929 30607 15963
rect 15485 15861 15519 15895
rect 19257 15861 19291 15895
rect 28733 15861 28767 15895
rect 31125 15861 31159 15895
rect 36829 15861 36863 15895
rect 37657 15861 37691 15895
rect 9873 15657 9907 15691
rect 17969 15589 18003 15623
rect 23213 15589 23247 15623
rect 30021 15589 30055 15623
rect 30573 15589 30607 15623
rect 2881 15521 2915 15555
rect 3433 15521 3467 15555
rect 9689 15521 9723 15555
rect 14933 15521 14967 15555
rect 22937 15521 22971 15555
rect 26709 15521 26743 15555
rect 27445 15521 27479 15555
rect 36461 15521 36495 15555
rect 36645 15521 36679 15555
rect 38301 15521 38335 15555
rect 4629 15453 4663 15487
rect 9597 15453 9631 15487
rect 12449 15453 12483 15487
rect 12633 15453 12667 15487
rect 12909 15453 12943 15487
rect 15200 15453 15234 15487
rect 17325 15453 17359 15487
rect 17509 15453 17543 15487
rect 17601 15453 17635 15487
rect 17693 15453 17727 15487
rect 19533 15453 19567 15487
rect 22845 15453 22879 15487
rect 27353 15453 27387 15487
rect 29009 15453 29043 15487
rect 29193 15453 29227 15487
rect 30202 15453 30236 15487
rect 30665 15453 30699 15487
rect 3249 15385 3283 15419
rect 4261 15385 4295 15419
rect 26464 15385 26498 15419
rect 29101 15385 29135 15419
rect 13093 15317 13127 15351
rect 16313 15317 16347 15351
rect 19625 15317 19659 15351
rect 25329 15317 25363 15351
rect 27721 15317 27755 15351
rect 30205 15317 30239 15351
rect 12909 15113 12943 15147
rect 20085 15113 20119 15147
rect 23581 15113 23615 15147
rect 26065 15113 26099 15147
rect 30665 15113 30699 15147
rect 24716 15045 24750 15079
rect 12449 14977 12483 15011
rect 12633 14977 12667 15011
rect 13369 14977 13403 15011
rect 13553 14977 13587 15011
rect 14105 14977 14139 15011
rect 14289 14977 14323 15011
rect 19257 14977 19291 15011
rect 19441 14977 19475 15011
rect 20026 14977 20060 15011
rect 21097 14977 21131 15011
rect 24961 14977 24995 15011
rect 25973 14977 26007 15011
rect 26157 14977 26191 15011
rect 30297 14977 30331 15011
rect 1869 14909 1903 14943
rect 2053 14909 2087 14943
rect 2789 14909 2823 14943
rect 12549 14909 12583 14943
rect 12725 14909 12759 14943
rect 20545 14909 20579 14943
rect 21281 14909 21315 14943
rect 30205 14909 30239 14943
rect 19901 14841 19935 14875
rect 20453 14841 20487 14875
rect 13461 14773 13495 14807
rect 14105 14773 14139 14807
rect 19441 14773 19475 14807
rect 1869 14569 1903 14603
rect 2697 14569 2731 14603
rect 16313 14569 16347 14603
rect 18245 14569 18279 14603
rect 19717 14569 19751 14603
rect 27261 14569 27295 14603
rect 27813 14569 27847 14603
rect 30021 14569 30055 14603
rect 22385 14501 22419 14535
rect 16129 14433 16163 14467
rect 16865 14433 16899 14467
rect 21097 14433 21131 14467
rect 2789 14365 2823 14399
rect 10333 14365 10367 14399
rect 15669 14365 15703 14399
rect 16405 14365 16439 14399
rect 20830 14365 20864 14399
rect 22109 14365 22143 14399
rect 27442 14365 27476 14399
rect 27905 14365 27939 14399
rect 10578 14297 10612 14331
rect 15402 14297 15436 14331
rect 17110 14297 17144 14331
rect 22385 14297 22419 14331
rect 29929 14297 29963 14331
rect 11713 14229 11747 14263
rect 14289 14229 14323 14263
rect 16129 14229 16163 14263
rect 22201 14229 22235 14263
rect 27445 14229 27479 14263
rect 2237 14025 2271 14059
rect 10241 14025 10275 14059
rect 12633 14025 12667 14059
rect 14197 14025 14231 14059
rect 14657 14025 14691 14059
rect 16221 14025 16255 14059
rect 18705 14025 18739 14059
rect 19809 14025 19843 14059
rect 20085 14025 20119 14059
rect 22109 14025 22143 14059
rect 25789 14025 25823 14059
rect 27905 14025 27939 14059
rect 14565 13957 14599 13991
rect 15393 13957 15427 13991
rect 19533 13957 19567 13991
rect 19901 13957 19935 13991
rect 21281 13957 21315 13991
rect 2329 13889 2363 13923
rect 10057 13889 10091 13923
rect 12725 13889 12759 13923
rect 15669 13889 15703 13923
rect 16129 13889 16163 13923
rect 16313 13889 16347 13923
rect 17141 13889 17175 13923
rect 18981 13889 19015 13923
rect 19073 13889 19107 13923
rect 19717 13889 19751 13923
rect 23222 13889 23256 13923
rect 23489 13889 23523 13923
rect 24409 13889 24443 13923
rect 24676 13889 24710 13923
rect 28273 13889 28307 13923
rect 29193 13889 29227 13923
rect 29377 13889 29411 13923
rect 29837 13889 29871 13923
rect 30113 13889 30147 13923
rect 14749 13821 14783 13855
rect 15393 13821 15427 13855
rect 16865 13821 16899 13855
rect 21465 13821 21499 13855
rect 28365 13821 28399 13855
rect 29009 13821 29043 13855
rect 15577 13753 15611 13787
rect 18889 13685 18923 13719
rect 9965 13481 9999 13515
rect 12633 13481 12667 13515
rect 13369 13481 13403 13515
rect 16957 13481 16991 13515
rect 17877 13481 17911 13515
rect 21925 13481 21959 13515
rect 22845 13481 22879 13515
rect 23765 13481 23799 13515
rect 25145 13481 25179 13515
rect 26709 13481 26743 13515
rect 17049 13413 17083 13447
rect 26157 13413 26191 13447
rect 10425 13345 10459 13379
rect 16865 13345 16899 13379
rect 13185 13277 13219 13311
rect 13369 13277 13403 13311
rect 17141 13277 17175 13311
rect 17601 13277 17635 13311
rect 22109 13277 22143 13311
rect 22293 13277 22327 13311
rect 22753 13277 22787 13311
rect 22937 13277 22971 13311
rect 24961 13277 24995 13311
rect 25145 13277 25179 13311
rect 26282 13277 26316 13311
rect 26801 13277 26835 13311
rect 27813 13277 27847 13311
rect 28089 13277 28123 13311
rect 37841 13277 37875 13311
rect 9597 13209 9631 13243
rect 9781 13209 9815 13243
rect 10692 13209 10726 13243
rect 12541 13209 12575 13243
rect 17785 13209 17819 13243
rect 23857 13209 23891 13243
rect 11805 13141 11839 13175
rect 26341 13141 26375 13175
rect 27629 13141 27663 13175
rect 27997 13141 28031 13175
rect 9505 12937 9539 12971
rect 10333 12937 10367 12971
rect 15393 12937 15427 12971
rect 17325 12937 17359 12971
rect 17969 12937 18003 12971
rect 26525 12937 26559 12971
rect 27813 12937 27847 12971
rect 10701 12869 10735 12903
rect 14749 12869 14783 12903
rect 15577 12869 15611 12903
rect 19533 12869 19567 12903
rect 2237 12801 2271 12835
rect 9137 12801 9171 12835
rect 10241 12801 10275 12835
rect 10609 12801 10643 12835
rect 13277 12801 13311 12835
rect 15301 12801 15335 12835
rect 16037 12801 16071 12835
rect 16221 12801 16255 12835
rect 17233 12801 17267 12835
rect 17417 12801 17451 12835
rect 18153 12801 18187 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 18521 12801 18555 12835
rect 19257 12801 19291 12835
rect 20177 12801 20211 12835
rect 20269 12801 20303 12835
rect 25145 12801 25179 12835
rect 26157 12801 26191 12835
rect 37473 12801 37507 12835
rect 9229 12733 9263 12767
rect 13001 12733 13035 12767
rect 19533 12733 19567 12767
rect 25237 12733 25271 12767
rect 26065 12733 26099 12767
rect 27353 12733 27387 12767
rect 28733 12733 28767 12767
rect 14565 12665 14599 12699
rect 15577 12665 15611 12699
rect 25513 12665 25547 12699
rect 27721 12665 27755 12699
rect 28365 12665 28399 12699
rect 2145 12597 2179 12631
rect 10517 12597 10551 12631
rect 12725 12597 12759 12631
rect 13185 12597 13219 12631
rect 16129 12597 16163 12631
rect 19349 12597 19383 12631
rect 19993 12597 20027 12631
rect 28273 12597 28307 12631
rect 37565 12597 37599 12631
rect 10609 12393 10643 12427
rect 13001 12393 13035 12427
rect 14473 12393 14507 12427
rect 16589 12393 16623 12427
rect 18245 12393 18279 12427
rect 19993 12393 20027 12427
rect 20453 12393 20487 12427
rect 21925 12393 21959 12427
rect 22109 12393 22143 12427
rect 28089 12393 28123 12427
rect 14565 12325 14599 12359
rect 15025 12325 15059 12359
rect 18797 12325 18831 12359
rect 21189 12325 21223 12359
rect 1777 12257 1811 12291
rect 2789 12257 2823 12291
rect 11621 12257 11655 12291
rect 11713 12257 11747 12291
rect 12541 12257 12575 12291
rect 12633 12257 12667 12291
rect 16313 12257 16347 12291
rect 37197 12257 37231 12291
rect 38117 12257 38151 12291
rect 38301 12257 38335 12291
rect 1593 12189 1627 12223
rect 10425 12189 10459 12223
rect 10609 12189 10643 12223
rect 11805 12189 11839 12223
rect 12817 12189 12851 12223
rect 14289 12189 14323 12223
rect 14657 12189 14691 12223
rect 14749 12189 14783 12223
rect 16129 12189 16163 12223
rect 16221 12189 16255 12223
rect 16405 12189 16439 12223
rect 17049 12189 17083 12223
rect 17233 12189 17267 12223
rect 17417 12189 17451 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 18705 12189 18739 12223
rect 18889 12189 18923 12223
rect 19901 12189 19935 12223
rect 20177 12189 20211 12223
rect 20269 12189 20303 12223
rect 20913 12189 20947 12223
rect 21741 12189 21775 12223
rect 21833 12189 21867 12223
rect 27905 12189 27939 12223
rect 28089 12189 28123 12223
rect 12081 12121 12115 12155
rect 21189 12121 21223 12155
rect 11989 12053 12023 12087
rect 21005 12053 21039 12087
rect 11989 11849 12023 11883
rect 14197 11849 14231 11883
rect 16313 11849 16347 11883
rect 22017 11849 22051 11883
rect 14933 11781 14967 11815
rect 15117 11781 15151 11815
rect 22169 11781 22203 11815
rect 22385 11781 22419 11815
rect 1869 11713 1903 11747
rect 9965 11713 9999 11747
rect 11805 11713 11839 11747
rect 12081 11713 12115 11747
rect 12817 11713 12851 11747
rect 14013 11713 14047 11747
rect 14289 11713 14323 11747
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 15945 11713 15979 11747
rect 16037 11713 16071 11747
rect 17049 11713 17083 11747
rect 18061 11713 18095 11747
rect 19809 11713 19843 11747
rect 20085 11713 20119 11747
rect 21189 11713 21223 11747
rect 21281 11713 21315 11747
rect 21465 11713 21499 11747
rect 37473 11713 37507 11747
rect 12725 11645 12759 11679
rect 13185 11645 13219 11679
rect 14749 11645 14783 11679
rect 16865 11645 16899 11679
rect 17325 11645 17359 11679
rect 18153 11645 18187 11679
rect 18429 11645 18463 11679
rect 19901 11645 19935 11679
rect 19993 11645 20027 11679
rect 20269 11645 20303 11679
rect 11805 11577 11839 11611
rect 13829 11577 13863 11611
rect 21465 11577 21499 11611
rect 10057 11509 10091 11543
rect 12541 11509 12575 11543
rect 17233 11509 17267 11543
rect 22201 11509 22235 11543
rect 37565 11509 37599 11543
rect 38301 11509 38335 11543
rect 12265 11305 12299 11339
rect 12633 11305 12667 11339
rect 14381 11305 14415 11339
rect 20361 11305 20395 11339
rect 16221 11237 16255 11271
rect 2973 11169 3007 11203
rect 9965 11169 9999 11203
rect 11621 11169 11655 11203
rect 11805 11169 11839 11203
rect 16037 11169 16071 11203
rect 37197 11169 37231 11203
rect 38117 11169 38151 11203
rect 38301 11169 38335 11203
rect 3433 11101 3467 11135
rect 12725 11101 12759 11135
rect 14473 11101 14507 11135
rect 16313 11101 16347 11135
rect 20269 11101 20303 11135
rect 20453 11101 20487 11135
rect 3249 11033 3283 11067
rect 16313 10965 16347 10999
rect 2789 10761 2823 10795
rect 2881 10625 2915 10659
rect 18429 10625 18463 10659
rect 2145 10557 2179 10591
rect 18613 10557 18647 10591
rect 19441 10557 19475 10591
rect 18521 10217 18555 10251
rect 18429 10013 18463 10047
rect 2513 9537 2547 9571
rect 23213 9537 23247 9571
rect 23857 9537 23891 9571
rect 23305 9469 23339 9503
rect 24041 9469 24075 9503
rect 25697 9469 25731 9503
rect 2053 9333 2087 9367
rect 2605 9333 2639 9367
rect 3249 8993 3283 9027
rect 3433 8993 3467 9027
rect 37841 8925 37875 8959
rect 1593 8857 1627 8891
rect 1869 8449 1903 8483
rect 1593 8381 1627 8415
rect 37841 8245 37875 8279
rect 37197 7905 37231 7939
rect 38301 7905 38335 7939
rect 38117 7769 38151 7803
rect 37565 7497 37599 7531
rect 37473 7361 37507 7395
rect 38117 7361 38151 7395
rect 2145 7157 2179 7191
rect 5365 7157 5399 7191
rect 38209 7157 38243 7191
rect 1593 6817 1627 6851
rect 3433 6817 3467 6851
rect 5365 6817 5399 6851
rect 5825 6817 5859 6851
rect 37197 6817 37231 6851
rect 38117 6817 38151 6851
rect 38301 6817 38335 6851
rect 3249 6681 3283 6715
rect 5549 6681 5583 6715
rect 2421 6409 2455 6443
rect 5549 6409 5583 6443
rect 2513 6273 2547 6307
rect 5457 6273 5491 6307
rect 37473 6273 37507 6307
rect 37565 6069 37599 6103
rect 37841 5729 37875 5763
rect 38117 5729 38151 5763
rect 1961 5661 1995 5695
rect 2789 5661 2823 5695
rect 3249 5661 3283 5695
rect 38301 5661 38335 5695
rect 3341 5525 3375 5559
rect 1869 5185 1903 5219
rect 37841 5185 37875 5219
rect 2053 5117 2087 5151
rect 2329 5117 2363 5151
rect 4169 4981 4203 5015
rect 36921 4981 36955 5015
rect 2237 4777 2271 4811
rect 37105 4641 37139 4675
rect 2329 4573 2363 4607
rect 2789 4573 2823 4607
rect 3985 4573 4019 4607
rect 4997 4573 5031 4607
rect 8309 4573 8343 4607
rect 25973 4573 26007 4607
rect 38209 4573 38243 4607
rect 38025 4505 38059 4539
rect 2881 4437 2915 4471
rect 5089 4437 5123 4471
rect 3801 4165 3835 4199
rect 8217 4097 8251 4131
rect 10517 4097 10551 4131
rect 24961 4097 24995 4131
rect 25973 4097 26007 4131
rect 37473 4097 37507 4131
rect 2973 4029 3007 4063
rect 3985 4029 4019 4063
rect 8401 4029 8435 4063
rect 8677 4029 8711 4063
rect 35817 4029 35851 4063
rect 36737 4029 36771 4063
rect 36921 4029 36955 4063
rect 38117 4029 38151 4063
rect 37565 3961 37599 3995
rect 4445 3893 4479 3927
rect 5549 3893 5583 3927
rect 10609 3893 10643 3927
rect 11805 3893 11839 3927
rect 19625 3893 19659 3927
rect 20729 3893 20763 3927
rect 22017 3893 22051 3927
rect 24869 3893 24903 3927
rect 26065 3893 26099 3927
rect 30021 3893 30055 3927
rect 33977 3893 34011 3927
rect 2789 3553 2823 3587
rect 3433 3553 3467 3587
rect 5549 3553 5583 3587
rect 5733 3553 5767 3587
rect 10609 3553 10643 3587
rect 10977 3553 11011 3587
rect 20729 3553 20763 3587
rect 21281 3553 21315 3587
rect 25881 3553 25915 3587
rect 26065 3553 26099 3587
rect 26433 3553 26467 3587
rect 30021 3553 30055 3587
rect 35909 3553 35943 3587
rect 4169 3485 4203 3519
rect 4997 3485 5031 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10425 3485 10459 3519
rect 13001 3485 13035 3519
rect 19625 3485 19659 3519
rect 19717 3485 19751 3519
rect 23213 3485 23247 3519
rect 24685 3485 24719 3519
rect 28365 3485 28399 3519
rect 29009 3485 29043 3519
rect 33885 3485 33919 3519
rect 35265 3485 35299 3519
rect 3249 3417 3283 3451
rect 7389 3417 7423 3451
rect 20913 3417 20947 3451
rect 29101 3417 29135 3451
rect 30205 3417 30239 3451
rect 31861 3417 31895 3451
rect 35357 3417 35391 3451
rect 36093 3417 36127 3451
rect 37749 3417 37783 3451
rect 4905 3349 4939 3383
rect 9229 3349 9263 3383
rect 28273 3349 28307 3383
rect 33977 3349 34011 3383
rect 37565 3145 37599 3179
rect 3525 3077 3559 3111
rect 4353 3077 4387 3111
rect 9045 3077 9079 3111
rect 19717 3077 19751 3111
rect 28089 3077 28123 3111
rect 34161 3077 34195 3111
rect 4169 3009 4203 3043
rect 8861 3009 8895 3043
rect 12265 3009 12299 3043
rect 12909 3009 12943 3043
rect 19533 3009 19567 3043
rect 22017 3009 22051 3043
rect 24317 3009 24351 3043
rect 33977 3009 34011 3043
rect 36277 3009 36311 3043
rect 37473 3009 37507 3043
rect 38117 3009 38151 3043
rect 2881 2941 2915 2975
rect 3709 2941 3743 2975
rect 4813 2941 4847 2975
rect 6561 2941 6595 2975
rect 6745 2941 6779 2975
rect 7757 2941 7791 2975
rect 9321 2941 9355 2975
rect 12357 2941 12391 2975
rect 13093 2941 13127 2975
rect 13553 2941 13587 2975
rect 19993 2941 20027 2975
rect 22201 2941 22235 2975
rect 22569 2941 22603 2975
rect 24501 2941 24535 2975
rect 24777 2941 24811 2975
rect 27905 2941 27939 2975
rect 28365 2941 28399 2975
rect 34805 2941 34839 2975
rect 2513 2601 2547 2635
rect 6745 2601 6779 2635
rect 7481 2601 7515 2635
rect 8493 2601 8527 2635
rect 9781 2601 9815 2635
rect 20821 2601 20855 2635
rect 22109 2601 22143 2635
rect 23029 2601 23063 2635
rect 27997 2601 28031 2635
rect 10333 2533 10367 2567
rect 31033 2533 31067 2567
rect 3985 2465 4019 2499
rect 4721 2465 4755 2499
rect 11805 2465 11839 2499
rect 12265 2465 12299 2499
rect 24593 2465 24627 2499
rect 24777 2465 24811 2499
rect 25145 2465 25179 2499
rect 30021 2465 30055 2499
rect 36461 2465 36495 2499
rect 36921 2465 36955 2499
rect 1685 2397 1719 2431
rect 2605 2397 2639 2431
rect 3249 2397 3283 2431
rect 7573 2397 7607 2431
rect 8585 2397 8619 2431
rect 9873 2397 9907 2431
rect 10517 2397 10551 2431
rect 10977 2397 11011 2431
rect 20729 2397 20763 2431
rect 22017 2397 22051 2431
rect 22937 2397 22971 2431
rect 29745 2397 29779 2431
rect 37565 2397 37599 2431
rect 1869 2329 1903 2363
rect 3341 2329 3375 2363
rect 4169 2329 4203 2363
rect 11069 2329 11103 2363
rect 11989 2329 12023 2363
rect 31217 2329 31251 2363
rect 36737 2329 36771 2363
rect 37657 2329 37691 2363
<< metal1 >>
rect 37826 37612 37832 37664
rect 37884 37652 37890 37664
rect 39298 37652 39304 37664
rect 37884 37624 39304 37652
rect 37884 37612 37890 37624
rect 39298 37612 39304 37624
rect 39356 37612 39362 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1857 37315 1915 37321
rect 1857 37281 1869 37315
rect 1903 37312 1915 37315
rect 2406 37312 2412 37324
rect 1903 37284 2412 37312
rect 1903 37281 1915 37284
rect 1857 37275 1915 37281
rect 2406 37272 2412 37284
rect 2464 37272 2470 37324
rect 18233 37315 18291 37321
rect 18233 37281 18245 37315
rect 18279 37312 18291 37315
rect 19150 37312 19156 37324
rect 18279 37284 19156 37312
rect 18279 37281 18291 37284
rect 18233 37275 18291 37281
rect 19150 37272 19156 37284
rect 19208 37272 19214 37324
rect 25774 37312 25780 37324
rect 25735 37284 25780 37312
rect 25774 37272 25780 37284
rect 25832 37272 25838 37324
rect 28626 37312 28632 37324
rect 28587 37284 28632 37312
rect 28626 37272 28632 37284
rect 28684 37272 28690 37324
rect 30282 37272 30288 37324
rect 30340 37312 30346 37324
rect 30377 37315 30435 37321
rect 30377 37312 30389 37315
rect 30340 37284 30389 37312
rect 30340 37272 30346 37284
rect 30377 37281 30389 37284
rect 30423 37281 30435 37315
rect 30377 37275 30435 37281
rect 32858 37272 32864 37324
rect 32916 37312 32922 37324
rect 32953 37315 33011 37321
rect 32953 37312 32965 37315
rect 32916 37284 32965 37312
rect 32916 37272 32922 37284
rect 32953 37281 32965 37284
rect 32999 37281 33011 37315
rect 32953 37275 33011 37281
rect 33042 37272 33048 37324
rect 33100 37312 33106 37324
rect 35342 37312 35348 37324
rect 33100 37284 35348 37312
rect 33100 37272 33106 37284
rect 35342 37272 35348 37284
rect 35400 37272 35406 37324
rect 38286 37312 38292 37324
rect 38247 37284 38292 37312
rect 38286 37272 38292 37284
rect 38344 37272 38350 37324
rect 14 37204 20 37256
rect 72 37244 78 37256
rect 1673 37247 1731 37253
rect 1673 37244 1685 37247
rect 72 37216 1685 37244
rect 72 37204 78 37216
rect 1673 37213 1685 37216
rect 1719 37213 1731 37247
rect 2498 37244 2504 37256
rect 2459 37216 2504 37244
rect 1673 37207 1731 37213
rect 2498 37204 2504 37216
rect 2556 37204 2562 37256
rect 3418 37244 3424 37256
rect 3379 37216 3424 37244
rect 3418 37204 3424 37216
rect 3476 37204 3482 37256
rect 4154 37244 4160 37256
rect 4115 37216 4160 37244
rect 4154 37204 4160 37216
rect 4212 37204 4218 37256
rect 4801 37247 4859 37253
rect 4801 37213 4813 37247
rect 4847 37213 4859 37247
rect 6546 37244 6552 37256
rect 6507 37216 6552 37244
rect 4801 37207 4859 37213
rect 4816 37176 4844 37207
rect 6546 37204 6552 37216
rect 6604 37204 6610 37256
rect 9214 37244 9220 37256
rect 9175 37216 9220 37244
rect 9214 37204 9220 37216
rect 9272 37204 9278 37256
rect 14458 37244 14464 37256
rect 14419 37216 14464 37244
rect 14458 37204 14464 37216
rect 14516 37204 14522 37256
rect 14918 37244 14924 37256
rect 14879 37216 14924 37244
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 15749 37247 15807 37253
rect 15749 37213 15761 37247
rect 15795 37244 15807 37247
rect 16206 37244 16212 37256
rect 15795 37216 16212 37244
rect 15795 37213 15807 37216
rect 15749 37207 15807 37213
rect 16206 37204 16212 37216
rect 16264 37244 16270 37256
rect 17586 37244 17592 37256
rect 16264 37216 17592 37244
rect 16264 37204 16270 37216
rect 17586 37204 17592 37216
rect 17644 37204 17650 37256
rect 18874 37244 18880 37256
rect 18835 37216 18880 37244
rect 18874 37204 18880 37216
rect 18932 37204 18938 37256
rect 19426 37204 19432 37256
rect 19484 37244 19490 37256
rect 19797 37247 19855 37253
rect 19797 37244 19809 37247
rect 19484 37216 19809 37244
rect 19484 37204 19490 37216
rect 19797 37213 19809 37216
rect 19843 37213 19855 37247
rect 20990 37244 20996 37256
rect 20951 37216 20996 37244
rect 19797 37207 19855 37213
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 22097 37247 22155 37253
rect 22097 37213 22109 37247
rect 22143 37213 22155 37247
rect 22738 37244 22744 37256
rect 22699 37216 22744 37244
rect 22097 37207 22155 37213
rect 5350 37176 5356 37188
rect 4816 37148 5356 37176
rect 5350 37136 5356 37148
rect 5408 37176 5414 37188
rect 22112 37176 22140 37207
rect 22738 37204 22744 37216
rect 22796 37204 22802 37256
rect 23566 37244 23572 37256
rect 23527 37216 23572 37244
rect 23566 37204 23572 37216
rect 23624 37204 23630 37256
rect 26605 37247 26663 37253
rect 26605 37213 26617 37247
rect 26651 37244 26663 37247
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 26651 37216 27169 37244
rect 26651 37213 26663 37216
rect 26605 37207 26663 37213
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27798 37244 27804 37256
rect 27759 37216 27804 37244
rect 27157 37207 27215 37213
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 29917 37247 29975 37253
rect 29917 37213 29929 37247
rect 29963 37213 29975 37247
rect 32490 37244 32496 37256
rect 32451 37216 32496 37244
rect 29917 37207 29975 37213
rect 26234 37176 26240 37188
rect 5408 37148 26240 37176
rect 5408 37136 5414 37148
rect 26234 37136 26240 37148
rect 26292 37136 26298 37188
rect 26418 37176 26424 37188
rect 26379 37148 26424 37176
rect 26418 37136 26424 37148
rect 26476 37136 26482 37188
rect 4338 37068 4344 37120
rect 4396 37108 4402 37120
rect 4709 37111 4767 37117
rect 4709 37108 4721 37111
rect 4396 37080 4721 37108
rect 4396 37068 4402 37080
rect 4709 37077 4721 37080
rect 4755 37077 4767 37111
rect 4709 37071 4767 37077
rect 14642 37068 14648 37120
rect 14700 37108 14706 37120
rect 15657 37111 15715 37117
rect 15657 37108 15669 37111
rect 14700 37080 15669 37108
rect 14700 37068 14706 37080
rect 15657 37077 15669 37080
rect 15703 37077 15715 37111
rect 15657 37071 15715 37077
rect 17497 37111 17555 37117
rect 17497 37077 17509 37111
rect 17543 37108 17555 37111
rect 18690 37108 18696 37120
rect 17543 37080 18696 37108
rect 17543 37077 17555 37080
rect 17497 37071 17555 37077
rect 18690 37068 18696 37080
rect 18748 37068 18754 37120
rect 22189 37111 22247 37117
rect 22189 37077 22201 37111
rect 22235 37108 22247 37111
rect 22278 37108 22284 37120
rect 22235 37080 22284 37108
rect 22235 37077 22247 37080
rect 22189 37071 22247 37077
rect 22278 37068 22284 37080
rect 22336 37068 22342 37120
rect 29932 37108 29960 37207
rect 32490 37204 32496 37216
rect 32548 37204 32554 37256
rect 36906 37204 36912 37256
rect 36964 37244 36970 37256
rect 38010 37244 38016 37256
rect 36964 37216 37009 37244
rect 37971 37216 38016 37244
rect 36964 37204 36970 37216
rect 38010 37204 38016 37216
rect 38068 37204 38074 37256
rect 30098 37176 30104 37188
rect 30059 37148 30104 37176
rect 30098 37136 30104 37148
rect 30156 37136 30162 37188
rect 32674 37176 32680 37188
rect 32635 37148 32680 37176
rect 32674 37136 32680 37148
rect 32732 37136 32738 37188
rect 35069 37179 35127 37185
rect 35069 37145 35081 37179
rect 35115 37176 35127 37179
rect 36725 37179 36783 37185
rect 35115 37148 35894 37176
rect 35115 37145 35127 37148
rect 35069 37139 35127 37145
rect 30650 37108 30656 37120
rect 29932 37080 30656 37108
rect 30650 37068 30656 37080
rect 30708 37068 30714 37120
rect 35866 37108 35894 37148
rect 36725 37145 36737 37179
rect 36771 37176 36783 37179
rect 38194 37176 38200 37188
rect 36771 37148 38200 37176
rect 36771 37145 36783 37148
rect 36725 37139 36783 37145
rect 38194 37136 38200 37148
rect 38252 37136 38258 37188
rect 38654 37108 38660 37120
rect 35866 37080 38660 37108
rect 38654 37068 38660 37080
rect 38712 37068 38718 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 17586 36864 17592 36916
rect 17644 36904 17650 36916
rect 23474 36904 23480 36916
rect 17644 36876 23480 36904
rect 17644 36864 17650 36876
rect 23474 36864 23480 36876
rect 23532 36864 23538 36916
rect 26234 36864 26240 36916
rect 26292 36904 26298 36916
rect 38194 36904 38200 36916
rect 26292 36876 35894 36904
rect 38155 36876 38200 36904
rect 26292 36864 26298 36876
rect 1854 36836 1860 36848
rect 1815 36808 1860 36836
rect 1854 36796 1860 36808
rect 1912 36796 1918 36848
rect 2498 36796 2504 36848
rect 2556 36836 2562 36848
rect 4338 36836 4344 36848
rect 2556 36808 3740 36836
rect 4299 36808 4344 36836
rect 2556 36796 2562 36808
rect 3712 36777 3740 36808
rect 4338 36796 4344 36808
rect 4396 36796 4402 36848
rect 14642 36836 14648 36848
rect 14603 36808 14648 36836
rect 14642 36796 14648 36808
rect 14700 36796 14706 36848
rect 16301 36839 16359 36845
rect 16301 36805 16313 36839
rect 16347 36836 16359 36839
rect 16758 36836 16764 36848
rect 16347 36808 16764 36836
rect 16347 36805 16359 36808
rect 16301 36799 16359 36805
rect 16758 36796 16764 36808
rect 16816 36796 16822 36848
rect 22278 36836 22284 36848
rect 22239 36808 22284 36836
rect 22278 36796 22284 36808
rect 22336 36796 22342 36848
rect 27798 36836 27804 36848
rect 27172 36808 27804 36836
rect 3697 36771 3755 36777
rect 3697 36737 3709 36771
rect 3743 36737 3755 36771
rect 4154 36768 4160 36780
rect 4115 36740 4160 36768
rect 3697 36731 3755 36737
rect 4154 36728 4160 36740
rect 4212 36728 4218 36780
rect 6546 36768 6552 36780
rect 6507 36740 6552 36768
rect 6546 36728 6552 36740
rect 6604 36728 6610 36780
rect 9214 36768 9220 36780
rect 9175 36740 9220 36768
rect 9214 36728 9220 36740
rect 9272 36728 9278 36780
rect 19150 36728 19156 36780
rect 19208 36768 19214 36780
rect 19208 36740 19253 36768
rect 19208 36728 19214 36740
rect 19426 36728 19432 36780
rect 19484 36768 19490 36780
rect 19613 36771 19671 36777
rect 19613 36768 19625 36771
rect 19484 36740 19625 36768
rect 19484 36728 19490 36740
rect 19613 36737 19625 36740
rect 19659 36737 19671 36771
rect 19613 36731 19671 36737
rect 23566 36728 23572 36780
rect 23624 36768 23630 36780
rect 27172 36777 27200 36808
rect 27798 36796 27804 36808
rect 27856 36796 27862 36848
rect 31754 36796 31760 36848
rect 31812 36836 31818 36848
rect 32493 36839 32551 36845
rect 32493 36836 32505 36839
rect 31812 36808 32505 36836
rect 31812 36796 31818 36808
rect 32493 36805 32505 36808
rect 32539 36805 32551 36839
rect 35866 36836 35894 36876
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 37458 36836 37464 36848
rect 35866 36808 37464 36836
rect 32493 36799 32551 36805
rect 37458 36796 37464 36808
rect 37516 36836 37522 36848
rect 37516 36808 38148 36836
rect 37516 36796 37522 36808
rect 38120 36777 38148 36808
rect 24397 36771 24455 36777
rect 24397 36768 24409 36771
rect 23624 36740 24409 36768
rect 23624 36728 23630 36740
rect 24397 36737 24409 36740
rect 24443 36737 24455 36771
rect 24397 36731 24455 36737
rect 27157 36771 27215 36777
rect 27157 36737 27169 36771
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 38105 36771 38163 36777
rect 38105 36737 38117 36771
rect 38151 36737 38163 36771
rect 38105 36731 38163 36737
rect 3510 36700 3516 36712
rect 3471 36672 3516 36700
rect 3510 36660 3516 36672
rect 3568 36660 3574 36712
rect 4617 36703 4675 36709
rect 4617 36669 4629 36703
rect 4663 36669 4675 36703
rect 4617 36663 4675 36669
rect 3234 36592 3240 36644
rect 3292 36632 3298 36644
rect 4632 36632 4660 36663
rect 6454 36660 6460 36712
rect 6512 36700 6518 36712
rect 6733 36703 6791 36709
rect 6733 36700 6745 36703
rect 6512 36672 6745 36700
rect 6512 36660 6518 36672
rect 6733 36669 6745 36672
rect 6779 36669 6791 36703
rect 7098 36700 7104 36712
rect 7059 36672 7104 36700
rect 6733 36663 6791 36669
rect 7098 36660 7104 36672
rect 7156 36660 7162 36712
rect 9398 36700 9404 36712
rect 9359 36672 9404 36700
rect 9398 36660 9404 36672
rect 9456 36660 9462 36712
rect 9674 36700 9680 36712
rect 9635 36672 9680 36700
rect 9674 36660 9680 36672
rect 9732 36660 9738 36712
rect 14461 36703 14519 36709
rect 14461 36669 14473 36703
rect 14507 36700 14519 36703
rect 14918 36700 14924 36712
rect 14507 36672 14924 36700
rect 14507 36669 14519 36672
rect 14461 36663 14519 36669
rect 14918 36660 14924 36672
rect 14976 36660 14982 36712
rect 18046 36700 18052 36712
rect 18007 36672 18052 36700
rect 18046 36660 18052 36672
rect 18104 36660 18110 36712
rect 18966 36700 18972 36712
rect 18927 36672 18972 36700
rect 18966 36660 18972 36672
rect 19024 36660 19030 36712
rect 19797 36703 19855 36709
rect 19797 36669 19809 36703
rect 19843 36700 19855 36703
rect 19886 36700 19892 36712
rect 19843 36672 19892 36700
rect 19843 36669 19855 36672
rect 19797 36663 19855 36669
rect 19886 36660 19892 36672
rect 19944 36660 19950 36712
rect 20622 36660 20628 36712
rect 20680 36700 20686 36712
rect 20717 36703 20775 36709
rect 20717 36700 20729 36703
rect 20680 36672 20729 36700
rect 20680 36660 20686 36672
rect 20717 36669 20729 36672
rect 20763 36669 20775 36703
rect 20717 36663 20775 36669
rect 22097 36703 22155 36709
rect 22097 36669 22109 36703
rect 22143 36700 22155 36703
rect 22738 36700 22744 36712
rect 22143 36672 22744 36700
rect 22143 36669 22155 36672
rect 22097 36663 22155 36669
rect 22738 36660 22744 36672
rect 22796 36660 22802 36712
rect 22830 36660 22836 36712
rect 22888 36700 22894 36712
rect 24578 36700 24584 36712
rect 22888 36672 22933 36700
rect 24539 36672 24584 36700
rect 22888 36660 22894 36672
rect 24578 36660 24584 36672
rect 24636 36660 24642 36712
rect 24857 36703 24915 36709
rect 24857 36669 24869 36703
rect 24903 36669 24915 36703
rect 27338 36700 27344 36712
rect 27299 36672 27344 36700
rect 24857 36663 24915 36669
rect 3292 36604 4660 36632
rect 3292 36592 3298 36604
rect 23842 36592 23848 36644
rect 23900 36632 23906 36644
rect 24872 36632 24900 36663
rect 27338 36660 27344 36672
rect 27396 36660 27402 36712
rect 27617 36703 27675 36709
rect 27617 36669 27629 36703
rect 27663 36669 27675 36703
rect 27617 36663 27675 36669
rect 29457 36703 29515 36709
rect 29457 36669 29469 36703
rect 29503 36669 29515 36703
rect 29638 36700 29644 36712
rect 29599 36672 29644 36700
rect 29457 36663 29515 36669
rect 23900 36604 24900 36632
rect 23900 36592 23906 36604
rect 26510 36592 26516 36644
rect 26568 36632 26574 36644
rect 27632 36632 27660 36663
rect 26568 36604 27660 36632
rect 26568 36592 26574 36604
rect 28442 36592 28448 36644
rect 28500 36632 28506 36644
rect 29472 36632 29500 36663
rect 29638 36660 29644 36672
rect 29696 36660 29702 36712
rect 29730 36660 29736 36712
rect 29788 36700 29794 36712
rect 29917 36703 29975 36709
rect 29917 36700 29929 36703
rect 29788 36672 29929 36700
rect 29788 36660 29794 36672
rect 29917 36669 29929 36672
rect 29963 36669 29975 36703
rect 32306 36700 32312 36712
rect 32267 36672 32312 36700
rect 29917 36663 29975 36669
rect 32306 36660 32312 36672
rect 32364 36660 32370 36712
rect 32769 36703 32827 36709
rect 32769 36669 32781 36703
rect 32815 36669 32827 36703
rect 34606 36700 34612 36712
rect 34567 36672 34612 36700
rect 32769 36663 32827 36669
rect 28500 36604 29500 36632
rect 28500 36592 28506 36604
rect 32214 36592 32220 36644
rect 32272 36632 32278 36644
rect 32784 36632 32812 36663
rect 34606 36660 34612 36672
rect 34664 36660 34670 36712
rect 34790 36700 34796 36712
rect 34751 36672 34796 36700
rect 34790 36660 34796 36672
rect 34848 36660 34854 36712
rect 34882 36660 34888 36712
rect 34940 36700 34946 36712
rect 35069 36703 35127 36709
rect 35069 36700 35081 36703
rect 34940 36672 35081 36700
rect 34940 36660 34946 36672
rect 35069 36669 35081 36672
rect 35115 36669 35127 36703
rect 35069 36663 35127 36669
rect 32272 36604 32812 36632
rect 32272 36592 32278 36604
rect 37182 36524 37188 36576
rect 37240 36564 37246 36576
rect 37461 36567 37519 36573
rect 37461 36564 37473 36567
rect 37240 36536 37473 36564
rect 37240 36524 37246 36536
rect 37461 36533 37473 36536
rect 37507 36533 37519 36567
rect 37461 36527 37519 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 6454 36360 6460 36372
rect 6415 36332 6460 36360
rect 6454 36320 6460 36332
rect 6512 36320 6518 36372
rect 9398 36360 9404 36372
rect 9359 36332 9404 36360
rect 9398 36320 9404 36332
rect 9456 36320 9462 36372
rect 19886 36360 19892 36372
rect 19847 36332 19892 36360
rect 19886 36320 19892 36332
rect 19944 36320 19950 36372
rect 23385 36363 23443 36369
rect 23385 36329 23397 36363
rect 23431 36360 23443 36363
rect 24578 36360 24584 36372
rect 23431 36332 24584 36360
rect 23431 36329 23443 36332
rect 23385 36323 23443 36329
rect 24578 36320 24584 36332
rect 24636 36320 24642 36372
rect 37366 36292 37372 36304
rect 36740 36264 37372 36292
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 3418 36184 3424 36236
rect 3476 36224 3482 36236
rect 3973 36227 4031 36233
rect 3973 36224 3985 36227
rect 3476 36196 3985 36224
rect 3476 36184 3482 36196
rect 3973 36193 3985 36196
rect 4019 36193 4031 36227
rect 3973 36187 4031 36193
rect 4154 36184 4160 36236
rect 4212 36224 4218 36236
rect 4433 36227 4491 36233
rect 4433 36224 4445 36227
rect 4212 36196 4445 36224
rect 4212 36184 4218 36196
rect 4433 36193 4445 36196
rect 4479 36193 4491 36227
rect 4433 36187 4491 36193
rect 14458 36184 14464 36236
rect 14516 36224 14522 36236
rect 14737 36227 14795 36233
rect 14737 36224 14749 36227
rect 14516 36196 14749 36224
rect 14516 36184 14522 36196
rect 14737 36193 14749 36196
rect 14783 36193 14795 36227
rect 16114 36224 16120 36236
rect 16075 36196 16120 36224
rect 14737 36187 14795 36193
rect 16114 36184 16120 36196
rect 16172 36184 16178 36236
rect 17402 36224 17408 36236
rect 17363 36196 17408 36224
rect 17402 36184 17408 36196
rect 17460 36184 17466 36236
rect 18690 36224 18696 36236
rect 18651 36196 18696 36224
rect 18690 36184 18696 36196
rect 18748 36184 18754 36236
rect 18874 36224 18880 36236
rect 18835 36196 18880 36224
rect 18874 36184 18880 36196
rect 18932 36184 18938 36236
rect 20990 36224 20996 36236
rect 20951 36196 20996 36224
rect 20990 36184 20996 36196
rect 21048 36184 21054 36236
rect 22094 36224 22100 36236
rect 22055 36196 22100 36224
rect 22094 36184 22100 36196
rect 22152 36184 22158 36236
rect 25130 36224 25136 36236
rect 25091 36196 25136 36224
rect 25130 36184 25136 36196
rect 25188 36184 25194 36236
rect 27062 36184 27068 36236
rect 27120 36224 27126 36236
rect 27341 36227 27399 36233
rect 27341 36224 27353 36227
rect 27120 36196 27353 36224
rect 27120 36184 27126 36196
rect 27341 36193 27353 36196
rect 27387 36193 27399 36227
rect 27341 36187 27399 36193
rect 28994 36184 29000 36236
rect 29052 36224 29058 36236
rect 30193 36227 30251 36233
rect 30193 36224 30205 36227
rect 29052 36196 30205 36224
rect 29052 36184 29058 36196
rect 30193 36193 30205 36196
rect 30239 36193 30251 36227
rect 30193 36187 30251 36193
rect 30926 36184 30932 36236
rect 30984 36224 30990 36236
rect 36740 36233 36768 36264
rect 37366 36252 37372 36264
rect 37424 36252 37430 36304
rect 32493 36227 32551 36233
rect 32493 36224 32505 36227
rect 30984 36196 32505 36224
rect 30984 36184 30990 36196
rect 32493 36193 32505 36196
rect 32539 36193 32551 36227
rect 32493 36187 32551 36193
rect 36725 36227 36783 36233
rect 36725 36193 36737 36227
rect 36771 36193 36783 36227
rect 37182 36224 37188 36236
rect 37143 36196 37188 36224
rect 36725 36187 36783 36193
rect 37182 36184 37188 36196
rect 37240 36184 37246 36236
rect 1578 36156 1584 36168
rect 1539 36128 1584 36156
rect 1578 36116 1584 36128
rect 1636 36116 1642 36168
rect 6362 36156 6368 36168
rect 6323 36128 6368 36156
rect 6362 36116 6368 36128
rect 6420 36116 6426 36168
rect 9309 36159 9367 36165
rect 9309 36125 9321 36159
rect 9355 36125 9367 36159
rect 9309 36119 9367 36125
rect 1762 36088 1768 36100
rect 1723 36060 1768 36088
rect 1762 36048 1768 36060
rect 1820 36048 1826 36100
rect 4154 36088 4160 36100
rect 4115 36060 4160 36088
rect 4154 36048 4160 36060
rect 4212 36048 4218 36100
rect 8478 35980 8484 36032
rect 8536 36020 8542 36032
rect 9324 36020 9352 36119
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 19981 36159 20039 36165
rect 19981 36156 19993 36159
rect 19392 36128 19993 36156
rect 19392 36116 19398 36128
rect 19981 36125 19993 36128
rect 20027 36125 20039 36159
rect 19981 36119 20039 36125
rect 23293 36159 23351 36165
rect 23293 36125 23305 36159
rect 23339 36125 23351 36159
rect 24578 36156 24584 36168
rect 24539 36128 24584 36156
rect 23293 36119 23351 36125
rect 14918 36088 14924 36100
rect 14879 36060 14924 36088
rect 14918 36048 14924 36060
rect 14976 36048 14982 36100
rect 21174 36088 21180 36100
rect 21135 36060 21180 36088
rect 21174 36048 21180 36060
rect 21232 36048 21238 36100
rect 23308 36032 23336 36119
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 26878 36156 26884 36168
rect 26839 36128 26884 36156
rect 26878 36116 26884 36128
rect 26936 36116 26942 36168
rect 29086 36116 29092 36168
rect 29144 36156 29150 36168
rect 29733 36159 29791 36165
rect 29733 36156 29745 36159
rect 29144 36128 29745 36156
rect 29144 36116 29150 36128
rect 29733 36125 29745 36128
rect 29779 36125 29791 36159
rect 32030 36156 32036 36168
rect 31991 36128 32036 36156
rect 29733 36119 29791 36125
rect 32030 36116 32036 36128
rect 32088 36116 32094 36168
rect 37642 36156 37648 36168
rect 37603 36128 37648 36156
rect 37642 36116 37648 36128
rect 37700 36116 37706 36168
rect 24762 36088 24768 36100
rect 24723 36060 24768 36088
rect 24762 36048 24768 36060
rect 24820 36048 24826 36100
rect 26602 36048 26608 36100
rect 26660 36088 26666 36100
rect 27065 36091 27123 36097
rect 27065 36088 27077 36091
rect 26660 36060 27077 36088
rect 26660 36048 26666 36060
rect 27065 36057 27077 36060
rect 27111 36057 27123 36091
rect 29914 36088 29920 36100
rect 29875 36060 29920 36088
rect 27065 36051 27123 36057
rect 29914 36048 29920 36060
rect 29972 36048 29978 36100
rect 32214 36088 32220 36100
rect 32175 36060 32220 36088
rect 32214 36048 32220 36060
rect 32272 36048 32278 36100
rect 37001 36091 37059 36097
rect 37001 36057 37013 36091
rect 37047 36088 37059 36091
rect 37737 36091 37795 36097
rect 37737 36088 37749 36091
rect 37047 36060 37749 36088
rect 37047 36057 37059 36060
rect 37001 36051 37059 36057
rect 37737 36057 37749 36060
rect 37783 36057 37795 36091
rect 37737 36051 37795 36057
rect 15194 36020 15200 36032
rect 8536 35992 15200 36020
rect 8536 35980 8542 35992
rect 15194 35980 15200 35992
rect 15252 35980 15258 36032
rect 23290 35980 23296 36032
rect 23348 36020 23354 36032
rect 25038 36020 25044 36032
rect 23348 35992 25044 36020
rect 23348 35980 23354 35992
rect 25038 35980 25044 35992
rect 25096 35980 25102 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1762 35776 1768 35828
rect 1820 35816 1826 35828
rect 2409 35819 2467 35825
rect 2409 35816 2421 35819
rect 1820 35788 2421 35816
rect 1820 35776 1826 35788
rect 2409 35785 2421 35788
rect 2455 35785 2467 35819
rect 2409 35779 2467 35785
rect 3053 35819 3111 35825
rect 3053 35785 3065 35819
rect 3099 35816 3111 35819
rect 3510 35816 3516 35828
rect 3099 35788 3516 35816
rect 3099 35785 3111 35788
rect 3053 35779 3111 35785
rect 3510 35776 3516 35788
rect 3568 35776 3574 35828
rect 3697 35819 3755 35825
rect 3697 35785 3709 35819
rect 3743 35816 3755 35819
rect 4154 35816 4160 35828
rect 3743 35788 4160 35816
rect 3743 35785 3755 35788
rect 3697 35779 3755 35785
rect 4154 35776 4160 35788
rect 4212 35776 4218 35828
rect 14918 35776 14924 35828
rect 14976 35816 14982 35828
rect 15105 35819 15163 35825
rect 15105 35816 15117 35819
rect 14976 35788 15117 35816
rect 14976 35776 14982 35788
rect 15105 35785 15117 35788
rect 15151 35785 15163 35819
rect 15105 35779 15163 35785
rect 15194 35776 15200 35828
rect 15252 35816 15258 35828
rect 18785 35819 18843 35825
rect 15252 35788 16574 35816
rect 15252 35776 15258 35788
rect 16546 35748 16574 35788
rect 18785 35785 18797 35819
rect 18831 35816 18843 35819
rect 18966 35816 18972 35828
rect 18831 35788 18972 35816
rect 18831 35785 18843 35788
rect 18785 35779 18843 35785
rect 18966 35776 18972 35788
rect 19024 35776 19030 35828
rect 21085 35819 21143 35825
rect 21085 35785 21097 35819
rect 21131 35816 21143 35819
rect 21174 35816 21180 35828
rect 21131 35788 21180 35816
rect 21131 35785 21143 35788
rect 21085 35779 21143 35785
rect 21174 35776 21180 35788
rect 21232 35776 21238 35828
rect 23661 35819 23719 35825
rect 23661 35785 23673 35819
rect 23707 35816 23719 35819
rect 24762 35816 24768 35828
rect 23707 35788 24768 35816
rect 23707 35785 23719 35788
rect 23661 35779 23719 35785
rect 24762 35776 24768 35788
rect 24820 35776 24826 35828
rect 25133 35819 25191 35825
rect 25133 35785 25145 35819
rect 25179 35816 25191 35819
rect 26418 35816 26424 35828
rect 25179 35788 26424 35816
rect 25179 35785 25191 35788
rect 25133 35779 25191 35785
rect 26418 35776 26424 35788
rect 26476 35776 26482 35828
rect 29914 35776 29920 35828
rect 29972 35816 29978 35828
rect 30009 35819 30067 35825
rect 30009 35816 30021 35819
rect 29972 35788 30021 35816
rect 29972 35776 29978 35788
rect 30009 35785 30021 35788
rect 30055 35785 30067 35819
rect 30009 35779 30067 35785
rect 30653 35819 30711 35825
rect 30653 35785 30665 35819
rect 30699 35816 30711 35819
rect 32214 35816 32220 35828
rect 30699 35788 32220 35816
rect 30699 35785 30711 35788
rect 30653 35779 30711 35785
rect 32214 35776 32220 35788
rect 32272 35776 32278 35828
rect 23290 35748 23296 35760
rect 16546 35720 23296 35748
rect 23290 35708 23296 35720
rect 23348 35708 23354 35760
rect 26053 35751 26111 35757
rect 26053 35717 26065 35751
rect 26099 35748 26111 35751
rect 27338 35748 27344 35760
rect 26099 35720 27344 35748
rect 26099 35717 26111 35720
rect 26053 35711 26111 35717
rect 27338 35708 27344 35720
rect 27396 35708 27402 35760
rect 27617 35751 27675 35757
rect 27617 35717 27629 35751
rect 27663 35748 27675 35751
rect 27706 35748 27712 35760
rect 27663 35720 27712 35748
rect 27663 35717 27675 35720
rect 27617 35711 27675 35717
rect 27706 35708 27712 35720
rect 27764 35708 27770 35760
rect 28626 35708 28632 35760
rect 28684 35748 28690 35760
rect 34425 35751 34483 35757
rect 28684 35720 29500 35748
rect 28684 35708 28690 35720
rect 1578 35640 1584 35692
rect 1636 35680 1642 35692
rect 1673 35683 1731 35689
rect 1673 35680 1685 35683
rect 1636 35652 1685 35680
rect 1636 35640 1642 35652
rect 1673 35649 1685 35652
rect 1719 35649 1731 35683
rect 1673 35643 1731 35649
rect 2501 35683 2559 35689
rect 2501 35649 2513 35683
rect 2547 35680 2559 35683
rect 2590 35680 2596 35692
rect 2547 35652 2596 35680
rect 2547 35649 2559 35652
rect 2501 35643 2559 35649
rect 2590 35640 2596 35652
rect 2648 35640 2654 35692
rect 3145 35683 3203 35689
rect 3145 35649 3157 35683
rect 3191 35680 3203 35683
rect 3326 35680 3332 35692
rect 3191 35652 3332 35680
rect 3191 35649 3203 35652
rect 3145 35643 3203 35649
rect 3326 35640 3332 35652
rect 3384 35640 3390 35692
rect 3605 35683 3663 35689
rect 3605 35649 3617 35683
rect 3651 35680 3663 35683
rect 3786 35680 3792 35692
rect 3651 35652 3792 35680
rect 3651 35649 3663 35652
rect 3605 35643 3663 35649
rect 3786 35640 3792 35652
rect 3844 35680 3850 35692
rect 6362 35680 6368 35692
rect 3844 35652 6368 35680
rect 3844 35640 3850 35652
rect 6362 35640 6368 35652
rect 6420 35640 6426 35692
rect 15194 35680 15200 35692
rect 15155 35652 15200 35680
rect 15194 35640 15200 35652
rect 15252 35640 15258 35692
rect 16942 35640 16948 35692
rect 17000 35680 17006 35692
rect 17109 35683 17167 35689
rect 17109 35680 17121 35683
rect 17000 35652 17121 35680
rect 17000 35640 17006 35652
rect 17109 35649 17121 35652
rect 17155 35649 17167 35683
rect 18874 35680 18880 35692
rect 18835 35652 18880 35680
rect 17109 35643 17167 35649
rect 18874 35640 18880 35652
rect 18932 35640 18938 35692
rect 20714 35640 20720 35692
rect 20772 35680 20778 35692
rect 20993 35683 21051 35689
rect 20993 35680 21005 35683
rect 20772 35652 21005 35680
rect 20772 35640 20778 35652
rect 20993 35649 21005 35652
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 23474 35640 23480 35692
rect 23532 35680 23538 35692
rect 23569 35683 23627 35689
rect 23569 35680 23581 35683
rect 23532 35652 23581 35680
rect 23532 35640 23538 35652
rect 23569 35649 23581 35652
rect 23615 35649 23627 35683
rect 23569 35643 23627 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35680 24455 35683
rect 24578 35680 24584 35692
rect 24443 35652 24584 35680
rect 24443 35649 24455 35652
rect 24397 35643 24455 35649
rect 24578 35640 24584 35652
rect 24636 35640 24642 35692
rect 25038 35680 25044 35692
rect 24999 35652 25044 35680
rect 25038 35640 25044 35652
rect 25096 35640 25102 35692
rect 25958 35680 25964 35692
rect 25919 35652 25964 35680
rect 25958 35640 25964 35652
rect 26016 35640 26022 35692
rect 29472 35689 29500 35720
rect 34425 35717 34437 35751
rect 34471 35748 34483 35751
rect 35342 35748 35348 35760
rect 34471 35720 35348 35748
rect 34471 35717 34483 35720
rect 34425 35711 34483 35717
rect 35342 35708 35348 35720
rect 35400 35708 35406 35760
rect 29457 35683 29515 35689
rect 29457 35649 29469 35683
rect 29503 35649 29515 35683
rect 29457 35643 29515 35649
rect 30101 35683 30159 35689
rect 30101 35649 30113 35683
rect 30147 35680 30159 35683
rect 30190 35680 30196 35692
rect 30147 35652 30196 35680
rect 30147 35649 30159 35652
rect 30101 35643 30159 35649
rect 30190 35640 30196 35652
rect 30248 35640 30254 35692
rect 30558 35680 30564 35692
rect 30519 35652 30564 35680
rect 30558 35640 30564 35652
rect 30616 35640 30622 35692
rect 31389 35683 31447 35689
rect 31389 35649 31401 35683
rect 31435 35680 31447 35683
rect 32030 35680 32036 35692
rect 31435 35652 32036 35680
rect 31435 35649 31447 35652
rect 31389 35643 31447 35649
rect 32030 35640 32036 35652
rect 32088 35640 32094 35692
rect 38105 35683 38163 35689
rect 38105 35649 38117 35683
rect 38151 35680 38163 35683
rect 38194 35680 38200 35692
rect 38151 35652 38200 35680
rect 38151 35649 38163 35652
rect 38105 35643 38163 35649
rect 38194 35640 38200 35652
rect 38252 35640 38258 35692
rect 15286 35572 15292 35624
rect 15344 35612 15350 35624
rect 16853 35615 16911 35621
rect 16853 35612 16865 35615
rect 15344 35584 16865 35612
rect 15344 35572 15350 35584
rect 16853 35581 16865 35584
rect 16899 35581 16911 35615
rect 16853 35575 16911 35581
rect 27982 35572 27988 35624
rect 28040 35612 28046 35624
rect 29273 35615 29331 35621
rect 29273 35612 29285 35615
rect 28040 35584 29285 35612
rect 28040 35572 28046 35584
rect 29273 35581 29285 35584
rect 29319 35581 29331 35615
rect 33042 35612 33048 35624
rect 33003 35584 33048 35612
rect 29273 35575 29331 35581
rect 33042 35572 33048 35584
rect 33100 35572 33106 35624
rect 34609 35615 34667 35621
rect 34609 35581 34621 35615
rect 34655 35612 34667 35615
rect 34698 35612 34704 35624
rect 34655 35584 34704 35612
rect 34655 35581 34667 35584
rect 34609 35575 34667 35581
rect 34698 35572 34704 35584
rect 34756 35572 34762 35624
rect 35713 35615 35771 35621
rect 35713 35581 35725 35615
rect 35759 35581 35771 35615
rect 35713 35575 35771 35581
rect 35728 35544 35756 35575
rect 35802 35572 35808 35624
rect 35860 35612 35866 35624
rect 36725 35615 36783 35621
rect 36725 35612 36737 35615
rect 35860 35584 36737 35612
rect 35860 35572 35866 35584
rect 36725 35581 36737 35584
rect 36771 35581 36783 35615
rect 36725 35575 36783 35581
rect 36909 35615 36967 35621
rect 36909 35581 36921 35615
rect 36955 35612 36967 35615
rect 37461 35615 37519 35621
rect 37461 35612 37473 35615
rect 36955 35584 37473 35612
rect 36955 35581 36967 35584
rect 36909 35575 36967 35581
rect 37461 35581 37473 35584
rect 37507 35581 37519 35615
rect 37461 35575 37519 35581
rect 37918 35544 37924 35556
rect 35728 35516 37924 35544
rect 37918 35504 37924 35516
rect 37976 35504 37982 35556
rect 17862 35436 17868 35488
rect 17920 35476 17926 35488
rect 18233 35479 18291 35485
rect 18233 35476 18245 35479
rect 17920 35448 18245 35476
rect 17920 35436 17926 35448
rect 18233 35445 18245 35448
rect 18279 35445 18291 35479
rect 18233 35439 18291 35445
rect 36722 35436 36728 35488
rect 36780 35476 36786 35488
rect 38197 35479 38255 35485
rect 38197 35476 38209 35479
rect 36780 35448 38209 35476
rect 36780 35436 36786 35448
rect 38197 35445 38209 35448
rect 38243 35445 38255 35479
rect 38197 35439 38255 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 16942 35272 16948 35284
rect 16903 35244 16948 35272
rect 16942 35232 16948 35244
rect 17000 35232 17006 35284
rect 18690 35272 18696 35284
rect 18651 35244 18696 35272
rect 18690 35232 18696 35244
rect 18748 35232 18754 35284
rect 18874 35232 18880 35284
rect 18932 35272 18938 35284
rect 26602 35272 26608 35284
rect 18932 35244 26234 35272
rect 26563 35244 26608 35272
rect 18932 35232 18938 35244
rect 15378 35164 15384 35216
rect 15436 35204 15442 35216
rect 18892 35204 18920 35232
rect 15436 35176 18920 35204
rect 26206 35204 26234 35244
rect 26602 35232 26608 35244
rect 26660 35232 26666 35284
rect 26878 35232 26884 35284
rect 26936 35272 26942 35284
rect 27157 35275 27215 35281
rect 27157 35272 27169 35275
rect 26936 35244 27169 35272
rect 26936 35232 26942 35244
rect 27157 35241 27169 35244
rect 27203 35241 27215 35275
rect 27982 35272 27988 35284
rect 27943 35244 27988 35272
rect 27157 35235 27215 35241
rect 27982 35232 27988 35244
rect 28040 35232 28046 35284
rect 28629 35275 28687 35281
rect 28629 35241 28641 35275
rect 28675 35272 28687 35275
rect 29638 35272 29644 35284
rect 28675 35244 29644 35272
rect 28675 35241 28687 35244
rect 28629 35235 28687 35241
rect 29638 35232 29644 35244
rect 29696 35232 29702 35284
rect 30098 35272 30104 35284
rect 30059 35244 30104 35272
rect 30098 35232 30104 35244
rect 30156 35232 30162 35284
rect 30650 35272 30656 35284
rect 30611 35244 30656 35272
rect 30650 35232 30656 35244
rect 30708 35232 30714 35284
rect 31754 35272 31760 35284
rect 31715 35244 31760 35272
rect 31754 35232 31760 35244
rect 31812 35232 31818 35284
rect 32306 35272 32312 35284
rect 32267 35244 32312 35272
rect 32306 35232 32312 35244
rect 32364 35232 32370 35284
rect 32674 35232 32680 35284
rect 32732 35272 32738 35284
rect 33045 35275 33103 35281
rect 33045 35272 33057 35275
rect 32732 35244 33057 35272
rect 32732 35232 32738 35244
rect 33045 35241 33057 35244
rect 33091 35241 33103 35275
rect 33045 35235 33103 35241
rect 34333 35275 34391 35281
rect 34333 35241 34345 35275
rect 34379 35272 34391 35275
rect 34606 35272 34612 35284
rect 34379 35244 34612 35272
rect 34379 35241 34391 35244
rect 34333 35235 34391 35241
rect 34606 35232 34612 35244
rect 34664 35232 34670 35284
rect 34790 35232 34796 35284
rect 34848 35272 34854 35284
rect 34977 35275 35035 35281
rect 34977 35272 34989 35275
rect 34848 35244 34989 35272
rect 34848 35232 34854 35244
rect 34977 35241 34989 35244
rect 35023 35241 35035 35275
rect 34977 35235 35035 35241
rect 35713 35275 35771 35281
rect 35713 35241 35725 35275
rect 35759 35272 35771 35275
rect 35802 35272 35808 35284
rect 35759 35244 35808 35272
rect 35759 35241 35771 35244
rect 35713 35235 35771 35241
rect 35802 35232 35808 35244
rect 35860 35232 35866 35284
rect 30190 35204 30196 35216
rect 26206 35176 28672 35204
rect 15436 35164 15442 35176
rect 19521 35139 19579 35145
rect 19521 35136 19533 35139
rect 18800 35108 19533 35136
rect 14277 35071 14335 35077
rect 14277 35037 14289 35071
rect 14323 35068 14335 35071
rect 15286 35068 15292 35080
rect 14323 35040 15292 35068
rect 14323 35037 14335 35040
rect 14277 35031 14335 35037
rect 15286 35028 15292 35040
rect 15344 35028 15350 35080
rect 17129 35071 17187 35077
rect 17129 35037 17141 35071
rect 17175 35068 17187 35071
rect 17586 35068 17592 35080
rect 17175 35040 17592 35068
rect 17175 35037 17187 35040
rect 17129 35031 17187 35037
rect 17586 35028 17592 35040
rect 17644 35028 17650 35080
rect 18800 35012 18828 35108
rect 19521 35105 19533 35108
rect 19567 35105 19579 35139
rect 19521 35099 19579 35105
rect 19628 35108 21404 35136
rect 19426 35028 19432 35080
rect 19484 35068 19490 35080
rect 19628 35077 19656 35108
rect 19613 35071 19671 35077
rect 19613 35068 19625 35071
rect 19484 35040 19625 35068
rect 19484 35028 19490 35040
rect 19613 35037 19625 35040
rect 19659 35037 19671 35071
rect 19613 35031 19671 35037
rect 20625 35071 20683 35077
rect 20625 35037 20637 35071
rect 20671 35068 20683 35071
rect 20990 35068 20996 35080
rect 20671 35040 20996 35068
rect 20671 35037 20683 35040
rect 20625 35031 20683 35037
rect 20990 35028 20996 35040
rect 21048 35028 21054 35080
rect 21266 35068 21272 35080
rect 21227 35040 21272 35068
rect 21266 35028 21272 35040
rect 21324 35028 21330 35080
rect 21376 35068 21404 35108
rect 25038 35096 25044 35148
rect 25096 35136 25102 35148
rect 25096 35108 28580 35136
rect 25096 35096 25102 35108
rect 23382 35068 23388 35080
rect 21376 35040 23388 35068
rect 23382 35028 23388 35040
rect 23440 35028 23446 35080
rect 26510 35068 26516 35080
rect 26471 35040 26516 35068
rect 26510 35028 26516 35040
rect 26568 35068 26574 35080
rect 28552 35077 28580 35108
rect 28077 35071 28135 35077
rect 28077 35068 28089 35071
rect 26568 35040 28089 35068
rect 26568 35028 26574 35040
rect 28077 35037 28089 35040
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 28537 35071 28595 35077
rect 28537 35037 28549 35071
rect 28583 35037 28595 35071
rect 28537 35031 28595 35037
rect 14544 35003 14602 35009
rect 14544 34969 14556 35003
rect 14590 35000 14602 35003
rect 14642 35000 14648 35012
rect 14590 34972 14648 35000
rect 14590 34969 14602 34972
rect 14544 34963 14602 34969
rect 14642 34960 14648 34972
rect 14700 34960 14706 35012
rect 18677 35003 18735 35009
rect 18677 34969 18689 35003
rect 18723 35000 18735 35003
rect 18782 35000 18788 35012
rect 18723 34972 18788 35000
rect 18723 34969 18735 34972
rect 18677 34963 18735 34969
rect 18782 34960 18788 34972
rect 18840 34960 18846 35012
rect 18874 34960 18880 35012
rect 18932 35000 18938 35012
rect 21514 35003 21572 35009
rect 21514 35000 21526 35003
rect 18932 34972 18977 35000
rect 20824 34972 21526 35000
rect 18932 34960 18938 34972
rect 15654 34932 15660 34944
rect 15615 34904 15660 34932
rect 15654 34892 15660 34904
rect 15712 34892 15718 34944
rect 18138 34892 18144 34944
rect 18196 34932 18202 34944
rect 18509 34935 18567 34941
rect 18509 34932 18521 34935
rect 18196 34904 18521 34932
rect 18196 34892 18202 34904
rect 18509 34901 18521 34904
rect 18555 34901 18567 34935
rect 19978 34932 19984 34944
rect 19939 34904 19984 34932
rect 18509 34895 18567 34901
rect 19978 34892 19984 34904
rect 20036 34892 20042 34944
rect 20824 34941 20852 34972
rect 21514 34969 21526 34972
rect 21560 34969 21572 35003
rect 28644 35000 28672 35176
rect 30024 35176 30196 35204
rect 30024 35077 30052 35176
rect 30190 35164 30196 35176
rect 30248 35204 30254 35216
rect 33686 35204 33692 35216
rect 30248 35176 33692 35204
rect 30248 35164 30254 35176
rect 33686 35164 33692 35176
rect 33744 35164 33750 35216
rect 38194 35204 38200 35216
rect 33796 35176 38200 35204
rect 30009 35071 30067 35077
rect 30009 35037 30021 35071
rect 30055 35037 30067 35071
rect 30009 35031 30067 35037
rect 31665 35071 31723 35077
rect 31665 35037 31677 35071
rect 31711 35070 31723 35071
rect 33137 35071 33195 35077
rect 31711 35068 31800 35070
rect 31711 35042 33088 35068
rect 31711 35037 31723 35042
rect 31772 35040 33088 35042
rect 31665 35031 31723 35037
rect 32306 35000 32312 35012
rect 28644 34972 32312 35000
rect 21514 34963 21572 34969
rect 32306 34960 32312 34972
rect 32364 34960 32370 35012
rect 33060 35000 33088 35040
rect 33137 35037 33149 35071
rect 33183 35068 33195 35071
rect 33594 35068 33600 35080
rect 33183 35040 33600 35068
rect 33183 35037 33195 35040
rect 33137 35031 33195 35037
rect 33594 35028 33600 35040
rect 33652 35028 33658 35080
rect 33796 35000 33824 35176
rect 38194 35164 38200 35176
rect 38252 35164 38258 35216
rect 37642 35136 37648 35148
rect 35084 35108 37648 35136
rect 35084 35077 35112 35108
rect 37642 35096 37648 35108
rect 37700 35096 37706 35148
rect 37826 35136 37832 35148
rect 37787 35108 37832 35136
rect 37826 35096 37832 35108
rect 37884 35096 37890 35148
rect 35069 35071 35127 35077
rect 35069 35037 35081 35071
rect 35115 35037 35127 35071
rect 35069 35031 35127 35037
rect 35621 35071 35679 35077
rect 35621 35037 35633 35071
rect 35667 35037 35679 35071
rect 35621 35031 35679 35037
rect 33060 34972 33824 35000
rect 20809 34935 20867 34941
rect 20809 34901 20821 34935
rect 20855 34901 20867 34935
rect 20809 34895 20867 34901
rect 22370 34892 22376 34944
rect 22428 34932 22434 34944
rect 22649 34935 22707 34941
rect 22649 34932 22661 34935
rect 22428 34904 22661 34932
rect 22428 34892 22434 34904
rect 22649 34901 22661 34904
rect 22695 34901 22707 34935
rect 22649 34895 22707 34901
rect 25406 34892 25412 34944
rect 25464 34932 25470 34944
rect 25958 34932 25964 34944
rect 25464 34904 25964 34932
rect 25464 34892 25470 34904
rect 25958 34892 25964 34904
rect 26016 34932 26022 34944
rect 35636 34932 35664 35031
rect 38286 35028 38292 35080
rect 38344 35068 38350 35080
rect 38344 35040 38389 35068
rect 38344 35028 38350 35040
rect 37274 35000 37280 35012
rect 35866 34972 37280 35000
rect 35866 34932 35894 34972
rect 37274 34960 37280 34972
rect 37332 34960 37338 35012
rect 37550 34960 37556 35012
rect 37608 35000 37614 35012
rect 38105 35003 38163 35009
rect 38105 35000 38117 35003
rect 37608 34972 38117 35000
rect 37608 34960 37614 34972
rect 38105 34969 38117 34972
rect 38151 34969 38163 35003
rect 38105 34963 38163 34969
rect 26016 34904 35894 34932
rect 26016 34892 26022 34904
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2590 34688 2596 34740
rect 2648 34728 2654 34740
rect 2648 34700 6914 34728
rect 2648 34688 2654 34700
rect 6886 34660 6914 34700
rect 14826 34688 14832 34740
rect 14884 34728 14890 34740
rect 15930 34728 15936 34740
rect 14884 34700 15936 34728
rect 14884 34688 14890 34700
rect 15930 34688 15936 34700
rect 15988 34688 15994 34740
rect 17586 34728 17592 34740
rect 17547 34700 17592 34728
rect 17586 34688 17592 34700
rect 17644 34688 17650 34740
rect 19334 34728 19340 34740
rect 17696 34700 19340 34728
rect 17696 34660 17724 34700
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 20990 34728 20996 34740
rect 20951 34700 20996 34728
rect 20990 34688 20996 34700
rect 21048 34688 21054 34740
rect 30558 34688 30564 34740
rect 30616 34728 30622 34740
rect 37550 34728 37556 34740
rect 30616 34700 37412 34728
rect 37511 34700 37556 34728
rect 30616 34688 30622 34700
rect 6886 34632 17724 34660
rect 17773 34663 17831 34669
rect 17773 34629 17785 34663
rect 17819 34660 17831 34663
rect 18414 34660 18420 34672
rect 17819 34632 18420 34660
rect 17819 34629 17831 34632
rect 17773 34623 17831 34629
rect 18414 34620 18420 34632
rect 18472 34620 18478 34672
rect 18874 34620 18880 34672
rect 18932 34660 18938 34672
rect 22370 34660 22376 34672
rect 18932 34632 22376 34660
rect 18932 34620 18938 34632
rect 22370 34620 22376 34632
rect 22428 34620 22434 34672
rect 36722 34660 36728 34672
rect 36683 34632 36728 34660
rect 36722 34620 36728 34632
rect 36780 34620 36786 34672
rect 37384 34660 37412 34700
rect 37550 34688 37556 34700
rect 37608 34688 37614 34740
rect 37918 34660 37924 34672
rect 37384 34632 37924 34660
rect 37918 34620 37924 34632
rect 37976 34620 37982 34672
rect 2406 34552 2412 34604
rect 2464 34592 2470 34604
rect 2501 34595 2559 34601
rect 2501 34592 2513 34595
rect 2464 34564 2513 34592
rect 2464 34552 2470 34564
rect 2501 34561 2513 34564
rect 2547 34592 2559 34595
rect 3142 34592 3148 34604
rect 2547 34564 3148 34592
rect 2547 34561 2559 34564
rect 2501 34555 2559 34561
rect 3142 34552 3148 34564
rect 3200 34552 3206 34604
rect 15378 34592 15384 34604
rect 6886 34564 15384 34592
rect 3326 34524 3332 34536
rect 3287 34496 3332 34524
rect 3326 34484 3332 34496
rect 3384 34524 3390 34536
rect 6886 34524 6914 34564
rect 15378 34552 15384 34564
rect 15436 34552 15442 34604
rect 18138 34592 18144 34604
rect 18099 34564 18144 34592
rect 18138 34552 18144 34564
rect 18196 34552 18202 34604
rect 18693 34595 18751 34601
rect 18693 34561 18705 34595
rect 18739 34561 18751 34595
rect 18693 34555 18751 34561
rect 3384 34496 6914 34524
rect 14921 34527 14979 34533
rect 3384 34484 3390 34496
rect 14921 34493 14933 34527
rect 14967 34524 14979 34527
rect 15102 34524 15108 34536
rect 14967 34496 15108 34524
rect 14967 34493 14979 34496
rect 14921 34487 14979 34493
rect 15102 34484 15108 34496
rect 15160 34484 15166 34536
rect 17402 34484 17408 34536
rect 17460 34524 17466 34536
rect 17862 34524 17868 34536
rect 17460 34496 17868 34524
rect 17460 34484 17466 34496
rect 17862 34484 17868 34496
rect 17920 34524 17926 34536
rect 18708 34524 18736 34555
rect 19978 34552 19984 34604
rect 20036 34592 20042 34604
rect 20809 34595 20867 34601
rect 20809 34592 20821 34595
rect 20036 34564 20821 34592
rect 20036 34552 20042 34564
rect 20809 34561 20821 34564
rect 20855 34561 20867 34595
rect 22922 34592 22928 34604
rect 22883 34564 22928 34592
rect 20809 34555 20867 34561
rect 22922 34552 22928 34564
rect 22980 34552 22986 34604
rect 33594 34552 33600 34604
rect 33652 34592 33658 34604
rect 33689 34595 33747 34601
rect 33689 34592 33701 34595
rect 33652 34564 33701 34592
rect 33652 34552 33658 34564
rect 33689 34561 33701 34564
rect 33735 34561 33747 34595
rect 37458 34592 37464 34604
rect 37419 34564 37464 34592
rect 33689 34555 33747 34561
rect 37458 34552 37464 34564
rect 37516 34552 37522 34604
rect 38286 34592 38292 34604
rect 38247 34564 38292 34592
rect 38286 34552 38292 34564
rect 38344 34552 38350 34604
rect 17920 34496 18736 34524
rect 17920 34484 17926 34496
rect 18966 34484 18972 34536
rect 19024 34524 19030 34536
rect 19889 34527 19947 34533
rect 19889 34524 19901 34527
rect 19024 34496 19901 34524
rect 19024 34484 19030 34496
rect 19889 34493 19901 34496
rect 19935 34524 19947 34527
rect 19935 34496 20024 34524
rect 19935 34493 19947 34496
rect 19889 34487 19947 34493
rect 14645 34459 14703 34465
rect 14645 34425 14657 34459
rect 14691 34456 14703 34459
rect 14734 34456 14740 34468
rect 14691 34428 14740 34456
rect 14691 34425 14703 34428
rect 14645 34419 14703 34425
rect 14734 34416 14740 34428
rect 14792 34416 14798 34468
rect 19996 34456 20024 34496
rect 20070 34484 20076 34536
rect 20128 34524 20134 34536
rect 20165 34527 20223 34533
rect 20165 34524 20177 34527
rect 20128 34496 20177 34524
rect 20128 34484 20134 34496
rect 20165 34493 20177 34496
rect 20211 34493 20223 34527
rect 20625 34527 20683 34533
rect 20625 34524 20637 34527
rect 20165 34487 20223 34493
rect 20272 34496 20637 34524
rect 20272 34456 20300 34496
rect 20625 34493 20637 34496
rect 20671 34493 20683 34527
rect 20625 34487 20683 34493
rect 23017 34527 23075 34533
rect 23017 34493 23029 34527
rect 23063 34524 23075 34527
rect 23569 34527 23627 34533
rect 23569 34524 23581 34527
rect 23063 34496 23581 34524
rect 23063 34493 23075 34496
rect 23017 34487 23075 34493
rect 23569 34493 23581 34496
rect 23615 34493 23627 34527
rect 23750 34524 23756 34536
rect 23711 34496 23756 34524
rect 23569 34487 23627 34493
rect 23750 34484 23756 34496
rect 23808 34484 23814 34536
rect 24486 34524 24492 34536
rect 24447 34496 24492 34524
rect 24486 34484 24492 34496
rect 24544 34484 24550 34536
rect 35710 34524 35716 34536
rect 35671 34496 35716 34524
rect 35710 34484 35716 34496
rect 35768 34484 35774 34536
rect 36909 34527 36967 34533
rect 36909 34493 36921 34527
rect 36955 34524 36967 34527
rect 37642 34524 37648 34536
rect 36955 34496 37648 34524
rect 36955 34493 36967 34496
rect 36909 34487 36967 34493
rect 37642 34484 37648 34496
rect 37700 34484 37706 34536
rect 28442 34456 28448 34468
rect 17788 34428 18920 34456
rect 19996 34428 20300 34456
rect 28403 34428 28448 34456
rect 14458 34388 14464 34400
rect 14419 34360 14464 34388
rect 14458 34348 14464 34360
rect 14516 34348 14522 34400
rect 17788 34397 17816 34428
rect 17773 34391 17831 34397
rect 17773 34357 17785 34391
rect 17819 34357 17831 34391
rect 17773 34351 17831 34357
rect 18690 34348 18696 34400
rect 18748 34388 18754 34400
rect 18785 34391 18843 34397
rect 18785 34388 18797 34391
rect 18748 34360 18797 34388
rect 18748 34348 18754 34360
rect 18785 34357 18797 34360
rect 18831 34357 18843 34391
rect 18892 34388 18920 34428
rect 28442 34416 28448 34428
rect 28500 34416 28506 34468
rect 29086 34456 29092 34468
rect 29047 34428 29092 34456
rect 29086 34416 29092 34428
rect 29144 34416 29150 34468
rect 32490 34416 32496 34468
rect 32548 34456 32554 34468
rect 32677 34459 32735 34465
rect 32677 34456 32689 34459
rect 32548 34428 32689 34456
rect 32548 34416 32554 34428
rect 32677 34425 32689 34428
rect 32723 34425 32735 34459
rect 32677 34419 32735 34425
rect 20162 34388 20168 34400
rect 18892 34360 20168 34388
rect 18785 34351 18843 34357
rect 20162 34348 20168 34360
rect 20220 34348 20226 34400
rect 33778 34388 33784 34400
rect 33739 34360 33784 34388
rect 33778 34348 33784 34360
rect 33836 34348 33842 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 14642 34184 14648 34196
rect 14603 34156 14648 34184
rect 14642 34144 14648 34156
rect 14700 34144 14706 34196
rect 17037 34187 17095 34193
rect 17037 34153 17049 34187
rect 17083 34184 17095 34187
rect 18138 34184 18144 34196
rect 17083 34156 18144 34184
rect 17083 34153 17095 34156
rect 17037 34147 17095 34153
rect 18138 34144 18144 34156
rect 18196 34144 18202 34196
rect 18414 34184 18420 34196
rect 18375 34156 18420 34184
rect 18414 34144 18420 34156
rect 18472 34144 18478 34196
rect 20162 34144 20168 34196
rect 20220 34184 20226 34196
rect 20349 34187 20407 34193
rect 20349 34184 20361 34187
rect 20220 34156 20361 34184
rect 20220 34144 20226 34156
rect 20349 34153 20361 34156
rect 20395 34153 20407 34187
rect 23382 34184 23388 34196
rect 23295 34156 23388 34184
rect 20349 34147 20407 34153
rect 23382 34144 23388 34156
rect 23440 34184 23446 34196
rect 23440 34156 26234 34184
rect 23440 34144 23446 34156
rect 15105 34051 15163 34057
rect 15105 34017 15117 34051
rect 15151 34048 15163 34051
rect 15654 34048 15660 34060
rect 15151 34020 15660 34048
rect 15151 34017 15163 34020
rect 15105 34011 15163 34017
rect 15654 34008 15660 34020
rect 15712 34008 15718 34060
rect 26206 34048 26234 34156
rect 34698 34144 34704 34196
rect 34756 34184 34762 34196
rect 35161 34187 35219 34193
rect 35161 34184 35173 34187
rect 34756 34156 35173 34184
rect 34756 34144 34762 34156
rect 35161 34153 35173 34156
rect 35207 34153 35219 34187
rect 35161 34147 35219 34153
rect 35989 34187 36047 34193
rect 35989 34153 36001 34187
rect 36035 34184 36047 34187
rect 36906 34184 36912 34196
rect 36035 34156 36912 34184
rect 36035 34153 36047 34156
rect 35989 34147 36047 34153
rect 36906 34144 36912 34156
rect 36964 34144 36970 34196
rect 26970 34048 26976 34060
rect 26206 34020 26976 34048
rect 26970 34008 26976 34020
rect 27028 34008 27034 34060
rect 32217 34051 32275 34057
rect 32217 34017 32229 34051
rect 32263 34048 32275 34051
rect 33870 34048 33876 34060
rect 32263 34020 33876 34048
rect 32263 34017 32275 34020
rect 32217 34011 32275 34017
rect 33870 34008 33876 34020
rect 33928 34008 33934 34060
rect 34057 34051 34115 34057
rect 34057 34017 34069 34051
rect 34103 34048 34115 34051
rect 35434 34048 35440 34060
rect 34103 34020 35440 34048
rect 34103 34017 34115 34020
rect 34057 34011 34115 34017
rect 35434 34008 35440 34020
rect 35492 34008 35498 34060
rect 38286 34048 38292 34060
rect 38247 34020 38292 34048
rect 38286 34008 38292 34020
rect 38344 34008 38350 34060
rect 1854 33940 1860 33992
rect 1912 33980 1918 33992
rect 1949 33983 2007 33989
rect 1949 33980 1961 33983
rect 1912 33952 1961 33980
rect 1912 33940 1918 33952
rect 1949 33949 1961 33952
rect 1995 33949 2007 33983
rect 1949 33943 2007 33949
rect 2777 33983 2835 33989
rect 2777 33949 2789 33983
rect 2823 33980 2835 33983
rect 3786 33980 3792 33992
rect 2823 33952 3792 33980
rect 2823 33949 2835 33952
rect 2777 33943 2835 33949
rect 3786 33940 3792 33952
rect 3844 33940 3850 33992
rect 14458 33980 14464 33992
rect 14419 33952 14464 33980
rect 14458 33940 14464 33952
rect 14516 33940 14522 33992
rect 15381 33983 15439 33989
rect 15381 33949 15393 33983
rect 15427 33949 15439 33983
rect 16850 33980 16856 33992
rect 16811 33952 16856 33980
rect 15381 33943 15439 33949
rect 15102 33872 15108 33924
rect 15160 33912 15166 33924
rect 15396 33912 15424 33943
rect 16850 33940 16856 33952
rect 16908 33940 16914 33992
rect 17129 33983 17187 33989
rect 17129 33949 17141 33983
rect 17175 33980 17187 33983
rect 17954 33980 17960 33992
rect 17175 33952 17960 33980
rect 17175 33949 17187 33952
rect 17129 33943 17187 33949
rect 17954 33940 17960 33952
rect 18012 33940 18018 33992
rect 18601 33983 18659 33989
rect 18601 33949 18613 33983
rect 18647 33980 18659 33983
rect 18690 33980 18696 33992
rect 18647 33952 18696 33980
rect 18647 33949 18659 33952
rect 18601 33943 18659 33949
rect 18690 33940 18696 33952
rect 18748 33940 18754 33992
rect 18782 33940 18788 33992
rect 18840 33980 18846 33992
rect 18877 33983 18935 33989
rect 18877 33980 18889 33983
rect 18840 33952 18889 33980
rect 18840 33940 18846 33952
rect 18877 33949 18889 33952
rect 18923 33980 18935 33983
rect 19242 33980 19248 33992
rect 18923 33952 19248 33980
rect 18923 33949 18935 33952
rect 18877 33943 18935 33949
rect 19242 33940 19248 33952
rect 19300 33980 19306 33992
rect 19981 33983 20039 33989
rect 19981 33980 19993 33983
rect 19300 33952 19993 33980
rect 19300 33940 19306 33952
rect 19981 33949 19993 33952
rect 20027 33949 20039 33983
rect 21450 33980 21456 33992
rect 21363 33952 21456 33980
rect 19981 33943 20039 33949
rect 21450 33940 21456 33952
rect 21508 33980 21514 33992
rect 21508 33952 21864 33980
rect 21508 33940 21514 33952
rect 15160 33884 15424 33912
rect 20349 33915 20407 33921
rect 15160 33872 15166 33884
rect 20349 33881 20361 33915
rect 20395 33912 20407 33915
rect 20990 33912 20996 33924
rect 20395 33884 20996 33912
rect 20395 33881 20407 33884
rect 20349 33875 20407 33881
rect 20990 33872 20996 33884
rect 21048 33872 21054 33924
rect 21266 33872 21272 33924
rect 21324 33912 21330 33924
rect 21698 33915 21756 33921
rect 21698 33912 21710 33915
rect 21324 33884 21710 33912
rect 21324 33872 21330 33884
rect 21698 33881 21710 33884
rect 21744 33881 21756 33915
rect 21836 33912 21864 33952
rect 22462 33940 22468 33992
rect 22520 33980 22526 33992
rect 23293 33983 23351 33989
rect 23293 33980 23305 33983
rect 22520 33952 23305 33980
rect 22520 33940 22526 33952
rect 23293 33949 23305 33952
rect 23339 33949 23351 33983
rect 25958 33980 25964 33992
rect 23293 33943 23351 33949
rect 23400 33952 25964 33980
rect 23400 33912 23428 33952
rect 25958 33940 25964 33952
rect 26016 33940 26022 33992
rect 26786 33940 26792 33992
rect 26844 33980 26850 33992
rect 27157 33983 27215 33989
rect 27157 33980 27169 33983
rect 26844 33952 27169 33980
rect 26844 33940 26850 33952
rect 27157 33949 27169 33952
rect 27203 33949 27215 33983
rect 27157 33943 27215 33949
rect 27246 33940 27252 33992
rect 27304 33980 27310 33992
rect 27801 33983 27859 33989
rect 27801 33980 27813 33983
rect 27304 33952 27813 33980
rect 27304 33940 27310 33952
rect 27801 33949 27813 33952
rect 27847 33949 27859 33983
rect 27801 33943 27859 33949
rect 27890 33940 27896 33992
rect 27948 33980 27954 33992
rect 27985 33983 28043 33989
rect 27985 33980 27997 33983
rect 27948 33952 27997 33980
rect 27948 33940 27954 33952
rect 27985 33949 27997 33952
rect 28031 33949 28043 33983
rect 36446 33980 36452 33992
rect 36407 33952 36452 33980
rect 27985 33943 28043 33949
rect 21836 33884 23428 33912
rect 21698 33875 21756 33881
rect 25498 33872 25504 33924
rect 25556 33912 25562 33924
rect 25694 33915 25752 33921
rect 25694 33912 25706 33915
rect 25556 33884 25706 33912
rect 25556 33872 25562 33884
rect 25694 33881 25706 33884
rect 25740 33881 25752 33915
rect 25694 33875 25752 33881
rect 27341 33915 27399 33921
rect 27341 33881 27353 33915
rect 27387 33912 27399 33915
rect 28000 33912 28028 33943
rect 36446 33940 36452 33952
rect 36504 33940 36510 33992
rect 32398 33912 32404 33924
rect 27387 33884 28028 33912
rect 32359 33884 32404 33912
rect 27387 33881 27399 33884
rect 27341 33875 27399 33881
rect 32398 33872 32404 33884
rect 32456 33872 32462 33924
rect 36633 33915 36691 33921
rect 36633 33881 36645 33915
rect 36679 33912 36691 33915
rect 36814 33912 36820 33924
rect 36679 33884 36820 33912
rect 36679 33881 36691 33884
rect 36633 33875 36691 33881
rect 36814 33872 36820 33884
rect 36872 33872 36878 33924
rect 2038 33804 2044 33856
rect 2096 33844 2102 33856
rect 2685 33847 2743 33853
rect 2685 33844 2697 33847
rect 2096 33816 2697 33844
rect 2096 33804 2102 33816
rect 2685 33813 2697 33816
rect 2731 33813 2743 33847
rect 2685 33807 2743 33813
rect 16574 33804 16580 33856
rect 16632 33844 16638 33856
rect 16669 33847 16727 33853
rect 16669 33844 16681 33847
rect 16632 33816 16681 33844
rect 16632 33804 16638 33816
rect 16669 33813 16681 33816
rect 16715 33813 16727 33847
rect 16669 33807 16727 33813
rect 18506 33804 18512 33856
rect 18564 33844 18570 33856
rect 18785 33847 18843 33853
rect 18785 33844 18797 33847
rect 18564 33816 18797 33844
rect 18564 33804 18570 33816
rect 18785 33813 18797 33816
rect 18831 33844 18843 33847
rect 18874 33844 18880 33856
rect 18831 33816 18880 33844
rect 18831 33813 18843 33816
rect 18785 33807 18843 33813
rect 18874 33804 18880 33816
rect 18932 33804 18938 33856
rect 20533 33847 20591 33853
rect 20533 33813 20545 33847
rect 20579 33844 20591 33847
rect 21082 33844 21088 33856
rect 20579 33816 21088 33844
rect 20579 33813 20591 33816
rect 20533 33807 20591 33813
rect 21082 33804 21088 33816
rect 21140 33804 21146 33856
rect 22830 33844 22836 33856
rect 22791 33816 22836 33844
rect 22830 33804 22836 33816
rect 22888 33804 22894 33856
rect 24581 33847 24639 33853
rect 24581 33813 24593 33847
rect 24627 33844 24639 33847
rect 24670 33844 24676 33856
rect 24627 33816 24676 33844
rect 24627 33813 24639 33816
rect 24581 33807 24639 33813
rect 24670 33804 24676 33816
rect 24728 33804 24734 33856
rect 27154 33804 27160 33856
rect 27212 33844 27218 33856
rect 27893 33847 27951 33853
rect 27893 33844 27905 33847
rect 27212 33816 27905 33844
rect 27212 33804 27218 33816
rect 27893 33813 27905 33816
rect 27939 33813 27951 33847
rect 27893 33807 27951 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 16850 33600 16856 33652
rect 16908 33640 16914 33652
rect 17129 33643 17187 33649
rect 17129 33640 17141 33643
rect 16908 33612 17141 33640
rect 16908 33600 16914 33612
rect 17129 33609 17141 33612
rect 17175 33609 17187 33643
rect 17129 33603 17187 33609
rect 19242 33600 19248 33652
rect 19300 33640 19306 33652
rect 19705 33643 19763 33649
rect 19705 33640 19717 33643
rect 19300 33612 19717 33640
rect 19300 33600 19306 33612
rect 19705 33609 19717 33612
rect 19751 33609 19763 33643
rect 21266 33640 21272 33652
rect 21227 33612 21272 33640
rect 19705 33603 19763 33609
rect 21266 33600 21272 33612
rect 21324 33600 21330 33652
rect 23750 33640 23756 33652
rect 23711 33612 23756 33640
rect 23750 33600 23756 33612
rect 23808 33600 23814 33652
rect 25498 33640 25504 33652
rect 25459 33612 25504 33640
rect 25498 33600 25504 33612
rect 25556 33600 25562 33652
rect 27246 33640 27252 33652
rect 27207 33612 27252 33640
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 32398 33640 32404 33652
rect 32359 33612 32404 33640
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 35342 33600 35348 33652
rect 35400 33640 35406 33652
rect 36173 33643 36231 33649
rect 36173 33640 36185 33643
rect 35400 33612 36185 33640
rect 35400 33600 35406 33612
rect 36173 33609 36185 33612
rect 36219 33609 36231 33643
rect 36814 33640 36820 33652
rect 36775 33612 36820 33640
rect 36173 33603 36231 33609
rect 36814 33600 36820 33612
rect 36872 33600 36878 33652
rect 2038 33572 2044 33584
rect 1999 33544 2044 33572
rect 2038 33532 2044 33544
rect 2096 33532 2102 33584
rect 17221 33575 17279 33581
rect 17221 33541 17233 33575
rect 17267 33572 17279 33575
rect 17954 33572 17960 33584
rect 17267 33544 17960 33572
rect 17267 33541 17279 33544
rect 17221 33535 17279 33541
rect 17954 33532 17960 33544
rect 18012 33572 18018 33584
rect 18598 33572 18604 33584
rect 18012 33544 18604 33572
rect 18012 33532 18018 33544
rect 18598 33532 18604 33544
rect 18656 33532 18662 33584
rect 24486 33572 24492 33584
rect 24447 33544 24492 33572
rect 24486 33532 24492 33544
rect 24544 33532 24550 33584
rect 24705 33575 24763 33581
rect 24705 33541 24717 33575
rect 24751 33572 24763 33575
rect 25590 33572 25596 33584
rect 24751 33544 25596 33572
rect 24751 33541 24763 33544
rect 24705 33535 24763 33541
rect 25590 33532 25596 33544
rect 25648 33532 25654 33584
rect 33778 33572 33784 33584
rect 33739 33544 33784 33572
rect 33778 33532 33784 33544
rect 33836 33532 33842 33584
rect 36446 33532 36452 33584
rect 36504 33572 36510 33584
rect 36504 33544 38148 33572
rect 36504 33532 36510 33544
rect 1854 33504 1860 33516
rect 1815 33476 1860 33504
rect 1854 33464 1860 33476
rect 1912 33464 1918 33516
rect 15010 33504 15016 33516
rect 14971 33476 15016 33504
rect 15010 33464 15016 33476
rect 15068 33464 15074 33516
rect 15102 33464 15108 33516
rect 15160 33504 15166 33516
rect 17313 33507 17371 33513
rect 15160 33476 15205 33504
rect 15160 33464 15166 33476
rect 17313 33473 17325 33507
rect 17359 33504 17371 33507
rect 18138 33504 18144 33516
rect 17359 33476 18144 33504
rect 17359 33473 17371 33476
rect 17313 33467 17371 33473
rect 18138 33464 18144 33476
rect 18196 33464 18202 33516
rect 19886 33504 19892 33516
rect 19847 33476 19892 33504
rect 19886 33464 19892 33476
rect 19944 33464 19950 33516
rect 19981 33507 20039 33513
rect 19981 33473 19993 33507
rect 20027 33473 20039 33507
rect 19981 33467 20039 33473
rect 2774 33436 2780 33448
rect 2735 33408 2780 33436
rect 2774 33396 2780 33408
rect 2832 33396 2838 33448
rect 14645 33439 14703 33445
rect 14645 33405 14657 33439
rect 14691 33436 14703 33439
rect 14734 33436 14740 33448
rect 14691 33408 14740 33436
rect 14691 33405 14703 33408
rect 14645 33399 14703 33405
rect 14734 33396 14740 33408
rect 14792 33436 14798 33448
rect 16853 33439 16911 33445
rect 16853 33436 16865 33439
rect 14792 33408 16865 33436
rect 14792 33396 14798 33408
rect 16853 33405 16865 33408
rect 16899 33436 16911 33439
rect 18046 33436 18052 33448
rect 16899 33408 18052 33436
rect 16899 33405 16911 33408
rect 16853 33399 16911 33405
rect 18046 33396 18052 33408
rect 18104 33436 18110 33448
rect 18966 33436 18972 33448
rect 18104 33408 18972 33436
rect 18104 33396 18110 33408
rect 18966 33396 18972 33408
rect 19024 33396 19030 33448
rect 19996 33312 20024 33467
rect 20070 33464 20076 33516
rect 20128 33508 20134 33516
rect 20128 33504 20208 33508
rect 21082 33504 21088 33516
rect 20128 33476 20221 33504
rect 21043 33476 21088 33504
rect 20128 33464 20134 33476
rect 20180 33436 20208 33476
rect 21082 33464 21088 33476
rect 21140 33464 21146 33516
rect 23658 33504 23664 33516
rect 23619 33476 23664 33504
rect 23658 33464 23664 33476
rect 23716 33464 23722 33516
rect 25317 33507 25375 33513
rect 25317 33504 25329 33507
rect 24872 33476 25329 33504
rect 21266 33436 21272 33448
rect 20180 33408 21272 33436
rect 21266 33396 21272 33408
rect 21324 33396 21330 33448
rect 20254 33368 20260 33380
rect 20215 33340 20260 33368
rect 20254 33328 20260 33340
rect 20312 33328 20318 33380
rect 23658 33328 23664 33380
rect 23716 33368 23722 33380
rect 24872 33377 24900 33476
rect 25317 33473 25329 33476
rect 25363 33473 25375 33507
rect 25317 33467 25375 33473
rect 26970 33464 26976 33516
rect 27028 33504 27034 33516
rect 27157 33507 27215 33513
rect 27157 33504 27169 33507
rect 27028 33476 27169 33504
rect 27028 33464 27034 33476
rect 27157 33473 27169 33476
rect 27203 33473 27215 33507
rect 27157 33467 27215 33473
rect 27341 33507 27399 33513
rect 27341 33473 27353 33507
rect 27387 33473 27399 33507
rect 27341 33467 27399 33473
rect 27893 33507 27951 33513
rect 27893 33473 27905 33507
rect 27939 33504 27951 33507
rect 27982 33504 27988 33516
rect 27939 33476 27988 33504
rect 27939 33473 27951 33476
rect 27893 33467 27951 33473
rect 26786 33396 26792 33448
rect 26844 33436 26850 33448
rect 27356 33436 27384 33467
rect 27982 33464 27988 33476
rect 28040 33464 28046 33516
rect 32306 33504 32312 33516
rect 32267 33476 32312 33504
rect 32306 33464 32312 33476
rect 32364 33464 32370 33516
rect 36265 33507 36323 33513
rect 36265 33473 36277 33507
rect 36311 33473 36323 33507
rect 36265 33467 36323 33473
rect 36909 33507 36967 33513
rect 36909 33473 36921 33507
rect 36955 33504 36967 33507
rect 37458 33504 37464 33516
rect 36955 33476 37464 33504
rect 36955 33473 36967 33476
rect 36909 33467 36967 33473
rect 26844 33408 27384 33436
rect 33597 33439 33655 33445
rect 26844 33396 26850 33408
rect 33597 33405 33609 33439
rect 33643 33436 33655 33439
rect 33870 33436 33876 33448
rect 33643 33408 33876 33436
rect 33643 33405 33655 33408
rect 33597 33399 33655 33405
rect 33870 33396 33876 33408
rect 33928 33396 33934 33448
rect 34514 33436 34520 33448
rect 34475 33408 34520 33436
rect 34514 33396 34520 33408
rect 34572 33396 34578 33448
rect 36280 33436 36308 33467
rect 37458 33464 37464 33476
rect 37516 33464 37522 33516
rect 38120 33513 38148 33544
rect 38105 33507 38163 33513
rect 38105 33473 38117 33507
rect 38151 33473 38163 33507
rect 38105 33467 38163 33473
rect 37366 33436 37372 33448
rect 36280 33408 37372 33436
rect 37366 33396 37372 33408
rect 37424 33396 37430 33448
rect 24857 33371 24915 33377
rect 23716 33340 24808 33368
rect 23716 33328 23722 33340
rect 14826 33300 14832 33312
rect 14787 33272 14832 33300
rect 14826 33260 14832 33272
rect 14884 33260 14890 33312
rect 19978 33300 19984 33312
rect 19891 33272 19984 33300
rect 19978 33260 19984 33272
rect 20036 33300 20042 33312
rect 20622 33300 20628 33312
rect 20036 33272 20628 33300
rect 20036 33260 20042 33272
rect 20622 33260 20628 33272
rect 20680 33300 20686 33312
rect 21358 33300 21364 33312
rect 20680 33272 21364 33300
rect 20680 33260 20686 33272
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 24578 33260 24584 33312
rect 24636 33300 24642 33312
rect 24673 33303 24731 33309
rect 24673 33300 24685 33303
rect 24636 33272 24685 33300
rect 24636 33260 24642 33272
rect 24673 33269 24685 33272
rect 24719 33269 24731 33303
rect 24780 33300 24808 33340
rect 24857 33337 24869 33371
rect 24903 33337 24915 33371
rect 36354 33368 36360 33380
rect 24857 33331 24915 33337
rect 26206 33340 36360 33368
rect 26206 33300 26234 33340
rect 36354 33328 36360 33340
rect 36412 33328 36418 33380
rect 24780 33272 26234 33300
rect 27985 33303 28043 33309
rect 24673 33263 24731 33269
rect 27985 33269 27997 33303
rect 28031 33300 28043 33303
rect 28166 33300 28172 33312
rect 28031 33272 28172 33300
rect 28031 33269 28043 33272
rect 27985 33263 28043 33269
rect 28166 33260 28172 33272
rect 28224 33260 28230 33312
rect 36446 33260 36452 33312
rect 36504 33300 36510 33312
rect 37461 33303 37519 33309
rect 37461 33300 37473 33303
rect 36504 33272 37473 33300
rect 36504 33260 36510 33272
rect 37461 33269 37473 33272
rect 37507 33269 37519 33303
rect 37461 33263 37519 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 20990 33096 20996 33108
rect 19306 33068 20576 33096
rect 20951 33068 20996 33096
rect 2225 32895 2283 32901
rect 2225 32861 2237 32895
rect 2271 32892 2283 32895
rect 3878 32892 3884 32904
rect 2271 32864 3884 32892
rect 2271 32861 2283 32864
rect 2225 32855 2283 32861
rect 3878 32852 3884 32864
rect 3936 32852 3942 32904
rect 10410 32892 10416 32904
rect 10371 32864 10416 32892
rect 10410 32852 10416 32864
rect 10468 32852 10474 32904
rect 10594 32892 10600 32904
rect 10555 32864 10600 32892
rect 10594 32852 10600 32864
rect 10652 32852 10658 32904
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32892 12955 32895
rect 14182 32892 14188 32904
rect 12943 32864 14188 32892
rect 12943 32861 12955 32864
rect 12897 32855 12955 32861
rect 14182 32852 14188 32864
rect 14240 32852 14246 32904
rect 14369 32895 14427 32901
rect 14369 32861 14381 32895
rect 14415 32892 14427 32895
rect 15194 32892 15200 32904
rect 14415 32864 15200 32892
rect 14415 32861 14427 32864
rect 14369 32855 14427 32861
rect 15194 32852 15200 32864
rect 15252 32852 15258 32904
rect 16301 32895 16359 32901
rect 16301 32861 16313 32895
rect 16347 32892 16359 32895
rect 18233 32895 18291 32901
rect 18233 32892 18245 32895
rect 16347 32864 16804 32892
rect 16347 32861 16359 32864
rect 16301 32855 16359 32861
rect 16776 32836 16804 32864
rect 17696 32864 18245 32892
rect 14642 32833 14648 32836
rect 14636 32787 14648 32833
rect 14700 32824 14706 32836
rect 16574 32833 16580 32836
rect 14700 32796 14736 32824
rect 14642 32784 14648 32787
rect 14700 32784 14706 32796
rect 16568 32787 16580 32833
rect 16632 32824 16638 32836
rect 16632 32796 16668 32824
rect 16574 32784 16580 32787
rect 16632 32784 16638 32796
rect 16758 32784 16764 32836
rect 16816 32784 16822 32836
rect 10502 32756 10508 32768
rect 10463 32728 10508 32756
rect 10502 32716 10508 32728
rect 10560 32716 10566 32768
rect 12710 32756 12716 32768
rect 12671 32728 12716 32756
rect 12710 32716 12716 32728
rect 12768 32716 12774 32768
rect 14918 32716 14924 32768
rect 14976 32756 14982 32768
rect 15749 32759 15807 32765
rect 15749 32756 15761 32759
rect 14976 32728 15761 32756
rect 14976 32716 14982 32728
rect 15749 32725 15761 32728
rect 15795 32725 15807 32759
rect 15749 32719 15807 32725
rect 17586 32716 17592 32768
rect 17644 32756 17650 32768
rect 17696 32765 17724 32864
rect 18233 32861 18245 32864
rect 18279 32861 18291 32895
rect 18233 32855 18291 32861
rect 18782 32852 18788 32904
rect 18840 32892 18846 32904
rect 19306 32892 19334 33068
rect 20070 32988 20076 33040
rect 20128 33028 20134 33040
rect 20128 33000 20300 33028
rect 20128 32988 20134 33000
rect 20272 32969 20300 33000
rect 20246 32963 20304 32969
rect 20246 32929 20258 32963
rect 20292 32929 20304 32963
rect 20246 32923 20304 32929
rect 18840 32864 19334 32892
rect 18840 32852 18846 32864
rect 19978 32852 19984 32904
rect 20036 32889 20042 32904
rect 20166 32895 20224 32901
rect 20166 32889 20178 32895
rect 20036 32861 20178 32889
rect 20212 32861 20224 32895
rect 20346 32892 20352 32904
rect 20307 32864 20352 32892
rect 20036 32852 20042 32861
rect 20166 32855 20224 32861
rect 20346 32852 20352 32864
rect 20404 32852 20410 32904
rect 20441 32895 20499 32901
rect 20441 32861 20453 32895
rect 20487 32892 20499 32895
rect 20548 32892 20576 33068
rect 20990 33056 20996 33068
rect 21048 33056 21054 33108
rect 26145 33099 26203 33105
rect 26145 33065 26157 33099
rect 26191 33096 26203 33099
rect 26789 33099 26847 33105
rect 26789 33096 26801 33099
rect 26191 33068 26801 33096
rect 26191 33065 26203 33068
rect 26145 33059 26203 33065
rect 26789 33065 26801 33068
rect 26835 33065 26847 33099
rect 26789 33059 26847 33065
rect 27062 33056 27068 33108
rect 27120 33096 27126 33108
rect 27120 33068 28396 33096
rect 27120 33056 27126 33068
rect 21358 32988 21364 33040
rect 21416 33028 21422 33040
rect 24857 33031 24915 33037
rect 21416 33000 23152 33028
rect 21416 32988 21422 33000
rect 21266 32920 21272 32972
rect 21324 32960 21330 32972
rect 21468 32969 21496 33000
rect 21453 32963 21511 32969
rect 21324 32932 21369 32960
rect 21324 32920 21330 32932
rect 21453 32929 21465 32963
rect 21499 32929 21511 32963
rect 21453 32923 21511 32929
rect 22281 32963 22339 32969
rect 22281 32929 22293 32963
rect 22327 32960 22339 32963
rect 22327 32932 22876 32960
rect 22327 32929 22339 32932
rect 22281 32923 22339 32929
rect 22848 32904 22876 32932
rect 21174 32892 21180 32904
rect 20487 32864 20576 32892
rect 21135 32864 21180 32892
rect 20487 32861 20499 32864
rect 20441 32855 20499 32861
rect 21174 32852 21180 32864
rect 21232 32852 21238 32904
rect 21358 32852 21364 32904
rect 21416 32892 21422 32904
rect 22370 32892 22376 32904
rect 21416 32864 21461 32892
rect 22331 32864 22376 32892
rect 21416 32852 21422 32864
rect 22370 32852 22376 32864
rect 22428 32852 22434 32904
rect 22830 32852 22836 32904
rect 22888 32892 22894 32904
rect 23124 32901 23152 33000
rect 24857 32997 24869 33031
rect 24903 33028 24915 33031
rect 24903 33000 25544 33028
rect 24903 32997 24915 33000
rect 24857 32991 24915 32997
rect 24946 32960 24952 32972
rect 24907 32932 24952 32960
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 25516 32960 25544 33000
rect 25590 32988 25596 33040
rect 25648 33028 25654 33040
rect 26329 33031 26387 33037
rect 26329 33028 26341 33031
rect 25648 33000 26341 33028
rect 25648 32988 25654 33000
rect 26329 32997 26341 33000
rect 26375 32997 26387 33031
rect 26329 32991 26387 32997
rect 26694 32988 26700 33040
rect 26752 33028 26758 33040
rect 26752 33000 27200 33028
rect 26752 32988 26758 33000
rect 26878 32960 26884 32972
rect 25516 32932 26884 32960
rect 26878 32920 26884 32932
rect 26936 32920 26942 32972
rect 22925 32895 22983 32901
rect 22925 32892 22937 32895
rect 22888 32864 22937 32892
rect 22888 32852 22894 32864
rect 22925 32861 22937 32864
rect 22971 32861 22983 32895
rect 22925 32855 22983 32861
rect 23109 32895 23167 32901
rect 23109 32861 23121 32895
rect 23155 32892 23167 32895
rect 26050 32892 26056 32904
rect 23155 32864 25820 32892
rect 26011 32864 26056 32892
rect 23155 32861 23167 32864
rect 23109 32855 23167 32861
rect 18417 32827 18475 32833
rect 18417 32793 18429 32827
rect 18463 32824 18475 32827
rect 18598 32824 18604 32836
rect 18463 32796 18604 32824
rect 18463 32793 18475 32796
rect 18417 32787 18475 32793
rect 18598 32784 18604 32796
rect 18656 32784 18662 32836
rect 18690 32784 18696 32836
rect 18748 32824 18754 32836
rect 22097 32827 22155 32833
rect 18748 32796 20116 32824
rect 18748 32784 18754 32796
rect 17681 32759 17739 32765
rect 17681 32756 17693 32759
rect 17644 32728 17693 32756
rect 17644 32716 17650 32728
rect 17681 32725 17693 32728
rect 17727 32725 17739 32759
rect 19978 32756 19984 32768
rect 19939 32728 19984 32756
rect 17681 32719 17739 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20088 32756 20116 32796
rect 22097 32793 22109 32827
rect 22143 32824 22155 32827
rect 22462 32824 22468 32836
rect 22143 32796 22468 32824
rect 22143 32793 22155 32796
rect 22097 32787 22155 32793
rect 22462 32784 22468 32796
rect 22520 32784 22526 32836
rect 24762 32824 24768 32836
rect 24723 32796 24768 32824
rect 24762 32784 24768 32796
rect 24820 32784 24826 32836
rect 25130 32824 25136 32836
rect 25091 32796 25136 32824
rect 25130 32784 25136 32796
rect 25188 32784 25194 32836
rect 25685 32827 25743 32833
rect 25685 32793 25697 32827
rect 25731 32793 25743 32827
rect 25792 32824 25820 32864
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 26145 32895 26203 32901
rect 26145 32861 26157 32895
rect 26191 32892 26203 32895
rect 26234 32892 26240 32904
rect 26191 32864 26240 32892
rect 26191 32861 26203 32864
rect 26145 32855 26203 32861
rect 26234 32852 26240 32864
rect 26292 32852 26298 32904
rect 26970 32852 26976 32904
rect 27028 32892 27034 32904
rect 27172 32901 27200 33000
rect 27356 33000 28120 33028
rect 27356 32904 27384 33000
rect 27065 32895 27123 32901
rect 27065 32892 27077 32895
rect 27028 32864 27077 32892
rect 27028 32852 27034 32864
rect 27065 32861 27077 32864
rect 27111 32861 27123 32895
rect 27065 32855 27123 32861
rect 27157 32895 27215 32901
rect 27157 32861 27169 32895
rect 27203 32861 27215 32895
rect 27157 32855 27215 32861
rect 27249 32895 27307 32901
rect 27249 32861 27261 32895
rect 27295 32892 27307 32895
rect 27338 32892 27344 32904
rect 27295 32864 27344 32892
rect 27295 32861 27307 32864
rect 27249 32855 27307 32861
rect 27338 32852 27344 32864
rect 27396 32852 27402 32904
rect 27430 32852 27436 32904
rect 27488 32892 27494 32904
rect 27890 32892 27896 32904
rect 27488 32864 27533 32892
rect 27851 32864 27896 32892
rect 27488 32852 27494 32864
rect 27890 32852 27896 32864
rect 27948 32852 27954 32904
rect 28092 32901 28120 33000
rect 28166 32920 28172 32972
rect 28224 32960 28230 32972
rect 28224 32932 28269 32960
rect 28224 32920 28230 32932
rect 28077 32895 28135 32901
rect 28077 32861 28089 32895
rect 28123 32861 28135 32895
rect 28258 32892 28264 32904
rect 28219 32864 28264 32892
rect 28077 32855 28135 32861
rect 28258 32852 28264 32864
rect 28316 32852 28322 32904
rect 28368 32901 28396 33068
rect 36446 32960 36452 32972
rect 36407 32932 36452 32960
rect 36446 32920 36452 32932
rect 36504 32920 36510 32972
rect 38286 32960 38292 32972
rect 38247 32932 38292 32960
rect 38286 32920 38292 32932
rect 38344 32920 38350 32972
rect 28353 32895 28411 32901
rect 28353 32861 28365 32895
rect 28399 32861 28411 32895
rect 28353 32855 28411 32861
rect 28994 32824 29000 32836
rect 25792 32796 29000 32824
rect 25685 32787 25743 32793
rect 22373 32759 22431 32765
rect 22373 32756 22385 32759
rect 20088 32728 22385 32756
rect 22373 32725 22385 32728
rect 22419 32725 22431 32759
rect 22373 32719 22431 32725
rect 25041 32759 25099 32765
rect 25041 32725 25053 32759
rect 25087 32756 25099 32759
rect 25700 32756 25728 32787
rect 28994 32784 29000 32796
rect 29052 32784 29058 32836
rect 36630 32824 36636 32836
rect 36591 32796 36636 32824
rect 36630 32784 36636 32796
rect 36688 32784 36694 32836
rect 25087 32728 25728 32756
rect 25087 32725 25099 32728
rect 25041 32719 25099 32725
rect 26602 32716 26608 32768
rect 26660 32756 26666 32768
rect 27154 32756 27160 32768
rect 26660 32728 27160 32756
rect 26660 32716 26666 32728
rect 27154 32716 27160 32728
rect 27212 32716 27218 32768
rect 27522 32716 27528 32768
rect 27580 32756 27586 32768
rect 28537 32759 28595 32765
rect 28537 32756 28549 32759
rect 27580 32728 28549 32756
rect 27580 32716 27586 32728
rect 28537 32725 28549 32728
rect 28583 32725 28595 32759
rect 28537 32719 28595 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 14642 32552 14648 32564
rect 14603 32524 14648 32552
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 24486 32512 24492 32564
rect 24544 32552 24550 32564
rect 24673 32555 24731 32561
rect 24673 32552 24685 32555
rect 24544 32524 24685 32552
rect 24544 32512 24550 32524
rect 24673 32521 24685 32524
rect 24719 32521 24731 32555
rect 24673 32515 24731 32521
rect 26050 32512 26056 32564
rect 26108 32552 26114 32564
rect 27525 32555 27583 32561
rect 27525 32552 27537 32555
rect 26108 32524 27537 32552
rect 26108 32512 26114 32524
rect 27525 32521 27537 32524
rect 27571 32521 27583 32555
rect 27525 32515 27583 32521
rect 36541 32555 36599 32561
rect 36541 32521 36553 32555
rect 36587 32552 36599 32555
rect 36630 32552 36636 32564
rect 36587 32524 36636 32552
rect 36587 32521 36599 32524
rect 36541 32515 36599 32521
rect 36630 32512 36636 32524
rect 36688 32512 36694 32564
rect 2498 32444 2504 32496
rect 2556 32484 2562 32496
rect 2556 32456 26740 32484
rect 2556 32444 2562 32456
rect 3878 32376 3884 32428
rect 3936 32416 3942 32428
rect 3936 32388 3981 32416
rect 3936 32376 3942 32388
rect 10502 32376 10508 32428
rect 10560 32416 10566 32428
rect 10882 32419 10940 32425
rect 10882 32416 10894 32419
rect 10560 32388 10894 32416
rect 10560 32376 10566 32388
rect 10882 32385 10894 32388
rect 10928 32385 10940 32419
rect 10882 32379 10940 32385
rect 12428 32419 12486 32425
rect 12428 32385 12440 32419
rect 12474 32416 12486 32419
rect 12710 32416 12716 32428
rect 12474 32388 12716 32416
rect 12474 32385 12486 32388
rect 12428 32379 12486 32385
rect 12710 32376 12716 32388
rect 12768 32376 12774 32428
rect 14826 32416 14832 32428
rect 14787 32388 14832 32416
rect 14826 32376 14832 32388
rect 14884 32376 14890 32428
rect 15010 32376 15016 32428
rect 15068 32416 15074 32428
rect 15105 32419 15163 32425
rect 15105 32416 15117 32419
rect 15068 32388 15117 32416
rect 15068 32376 15074 32388
rect 15105 32385 15117 32388
rect 15151 32416 15163 32419
rect 16022 32416 16028 32428
rect 15151 32388 16028 32416
rect 15151 32385 15163 32388
rect 15105 32379 15163 32385
rect 16022 32376 16028 32388
rect 16080 32376 16086 32428
rect 17402 32416 17408 32428
rect 17363 32388 17408 32416
rect 17402 32376 17408 32388
rect 17460 32376 17466 32428
rect 17586 32416 17592 32428
rect 17547 32388 17592 32416
rect 17586 32376 17592 32388
rect 17644 32416 17650 32428
rect 18233 32419 18291 32425
rect 18233 32416 18245 32419
rect 17644 32388 18245 32416
rect 17644 32376 17650 32388
rect 18233 32385 18245 32388
rect 18279 32385 18291 32419
rect 18506 32416 18512 32428
rect 18467 32388 18512 32416
rect 18233 32379 18291 32385
rect 18506 32376 18512 32388
rect 18564 32376 18570 32428
rect 18598 32376 18604 32428
rect 18656 32416 18662 32428
rect 19426 32416 19432 32428
rect 18656 32388 19288 32416
rect 19387 32388 19432 32416
rect 18656 32376 18662 32388
rect 2682 32348 2688 32360
rect 2643 32320 2688 32348
rect 2682 32308 2688 32320
rect 2740 32308 2746 32360
rect 3694 32348 3700 32360
rect 3655 32320 3700 32348
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 8665 32351 8723 32357
rect 8665 32317 8677 32351
rect 8711 32348 8723 32351
rect 8938 32348 8944 32360
rect 8711 32320 8944 32348
rect 8711 32317 8723 32320
rect 8665 32311 8723 32317
rect 8938 32308 8944 32320
rect 8996 32348 9002 32360
rect 11149 32351 11207 32357
rect 8996 32320 9812 32348
rect 8996 32308 9002 32320
rect 9033 32283 9091 32289
rect 9033 32249 9045 32283
rect 9079 32280 9091 32283
rect 9398 32280 9404 32292
rect 9079 32252 9404 32280
rect 9079 32249 9091 32252
rect 9033 32243 9091 32249
rect 9398 32240 9404 32252
rect 9456 32240 9462 32292
rect 9784 32289 9812 32320
rect 11149 32317 11161 32351
rect 11195 32348 11207 32351
rect 12158 32348 12164 32360
rect 11195 32320 12164 32348
rect 11195 32317 11207 32320
rect 11149 32311 11207 32317
rect 12158 32308 12164 32320
rect 12216 32308 12222 32360
rect 18049 32351 18107 32357
rect 18049 32317 18061 32351
rect 18095 32348 18107 32351
rect 19150 32348 19156 32360
rect 18095 32320 19156 32348
rect 18095 32317 18107 32320
rect 18049 32311 18107 32317
rect 19150 32308 19156 32320
rect 19208 32308 19214 32360
rect 19260 32348 19288 32388
rect 19426 32376 19432 32388
rect 19484 32376 19490 32428
rect 19889 32419 19947 32425
rect 19889 32416 19901 32419
rect 19536 32388 19901 32416
rect 19536 32348 19564 32388
rect 19889 32385 19901 32388
rect 19935 32416 19947 32419
rect 20806 32416 20812 32428
rect 19935 32388 20812 32416
rect 19935 32385 19947 32388
rect 19889 32379 19947 32385
rect 20806 32376 20812 32388
rect 20864 32376 20870 32428
rect 24670 32376 24676 32428
rect 24728 32416 24734 32428
rect 24857 32419 24915 32425
rect 24857 32416 24869 32419
rect 24728 32388 24869 32416
rect 24728 32376 24734 32388
rect 24857 32385 24869 32388
rect 24903 32385 24915 32419
rect 24857 32379 24915 32385
rect 25087 32419 25145 32425
rect 25087 32385 25099 32419
rect 25133 32416 25145 32419
rect 26602 32416 26608 32428
rect 25133 32388 26608 32416
rect 25133 32385 25145 32388
rect 25087 32379 25145 32385
rect 26602 32376 26608 32388
rect 26660 32376 26666 32428
rect 19260 32320 19564 32348
rect 19613 32351 19671 32357
rect 19613 32317 19625 32351
rect 19659 32348 19671 32351
rect 19978 32348 19984 32360
rect 19659 32320 19984 32348
rect 19659 32317 19671 32320
rect 19613 32311 19671 32317
rect 19978 32308 19984 32320
rect 20036 32308 20042 32360
rect 20254 32308 20260 32360
rect 20312 32348 20318 32360
rect 21177 32351 21235 32357
rect 21177 32348 21189 32351
rect 20312 32320 21189 32348
rect 20312 32308 20318 32320
rect 21177 32317 21189 32320
rect 21223 32348 21235 32351
rect 21358 32348 21364 32360
rect 21223 32320 21364 32348
rect 21223 32317 21235 32320
rect 21177 32311 21235 32317
rect 21358 32308 21364 32320
rect 21416 32308 21422 32360
rect 21453 32351 21511 32357
rect 21453 32317 21465 32351
rect 21499 32348 21511 32351
rect 22462 32348 22468 32360
rect 21499 32320 22468 32348
rect 21499 32317 21511 32320
rect 21453 32311 21511 32317
rect 9769 32283 9827 32289
rect 9769 32249 9781 32283
rect 9815 32249 9827 32283
rect 19245 32283 19303 32289
rect 19245 32280 19257 32283
rect 9769 32243 9827 32249
rect 13096 32252 19257 32280
rect 9125 32215 9183 32221
rect 9125 32181 9137 32215
rect 9171 32212 9183 32215
rect 9674 32212 9680 32224
rect 9171 32184 9680 32212
rect 9171 32181 9183 32184
rect 9125 32175 9183 32181
rect 9674 32172 9680 32184
rect 9732 32172 9738 32224
rect 9950 32172 9956 32224
rect 10008 32212 10014 32224
rect 13096 32212 13124 32252
rect 19245 32249 19257 32252
rect 19291 32249 19303 32283
rect 19245 32243 19303 32249
rect 20530 32240 20536 32292
rect 20588 32280 20594 32292
rect 21468 32280 21496 32311
rect 22462 32308 22468 32320
rect 22520 32308 22526 32360
rect 24949 32351 25007 32357
rect 24949 32317 24961 32351
rect 24995 32317 25007 32351
rect 25222 32348 25228 32360
rect 25183 32320 25228 32348
rect 24949 32311 25007 32317
rect 20588 32252 21496 32280
rect 20588 32240 20594 32252
rect 13538 32212 13544 32224
rect 10008 32184 13124 32212
rect 13499 32184 13544 32212
rect 10008 32172 10014 32184
rect 13538 32172 13544 32184
rect 13596 32172 13602 32224
rect 15013 32215 15071 32221
rect 15013 32181 15025 32215
rect 15059 32212 15071 32215
rect 15102 32212 15108 32224
rect 15059 32184 15108 32212
rect 15059 32181 15071 32184
rect 15013 32175 15071 32181
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 17221 32215 17279 32221
rect 17221 32181 17233 32215
rect 17267 32212 17279 32215
rect 17310 32212 17316 32224
rect 17267 32184 17316 32212
rect 17267 32181 17279 32184
rect 17221 32175 17279 32181
rect 17310 32172 17316 32184
rect 17368 32172 17374 32224
rect 18417 32215 18475 32221
rect 18417 32181 18429 32215
rect 18463 32212 18475 32215
rect 18782 32212 18788 32224
rect 18463 32184 18788 32212
rect 18463 32181 18475 32184
rect 18417 32175 18475 32181
rect 18782 32172 18788 32184
rect 18840 32172 18846 32224
rect 19610 32212 19616 32224
rect 19571 32184 19616 32212
rect 19610 32172 19616 32184
rect 19668 32172 19674 32224
rect 24964 32212 24992 32311
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 25314 32308 25320 32360
rect 25372 32348 25378 32360
rect 25372 32320 25417 32348
rect 25372 32308 25378 32320
rect 25498 32240 25504 32292
rect 25556 32280 25562 32292
rect 26712 32280 26740 32456
rect 26878 32444 26884 32496
rect 26936 32484 26942 32496
rect 28534 32484 28540 32496
rect 26936 32456 28540 32484
rect 26936 32444 26942 32456
rect 28534 32444 28540 32456
rect 28592 32444 28598 32496
rect 30558 32484 30564 32496
rect 28828 32456 30564 32484
rect 27154 32416 27160 32428
rect 27115 32388 27160 32416
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 27246 32376 27252 32428
rect 27304 32416 27310 32428
rect 27522 32416 27528 32428
rect 27304 32388 27349 32416
rect 27483 32388 27528 32416
rect 27304 32376 27310 32388
rect 27522 32376 27528 32388
rect 27580 32376 27586 32428
rect 28828 32416 28856 32456
rect 30558 32444 30564 32456
rect 30616 32444 30622 32496
rect 28994 32416 29000 32428
rect 27908 32388 28856 32416
rect 28955 32388 29000 32416
rect 27062 32308 27068 32360
rect 27120 32348 27126 32360
rect 27433 32351 27491 32357
rect 27433 32348 27445 32351
rect 27120 32320 27445 32348
rect 27120 32308 27126 32320
rect 27433 32317 27445 32320
rect 27479 32317 27491 32351
rect 27433 32311 27491 32317
rect 27908 32280 27936 32388
rect 28994 32376 29000 32388
rect 29052 32376 29058 32428
rect 36446 32416 36452 32428
rect 36407 32388 36452 32416
rect 36446 32376 36452 32388
rect 36504 32376 36510 32428
rect 37642 32416 37648 32428
rect 37603 32388 37648 32416
rect 37642 32376 37648 32388
rect 37700 32376 37706 32428
rect 29086 32348 29092 32360
rect 29047 32320 29092 32348
rect 29086 32308 29092 32320
rect 29144 32308 29150 32360
rect 25556 32252 26234 32280
rect 26712 32252 27936 32280
rect 25556 32240 25562 32252
rect 25038 32212 25044 32224
rect 24964 32184 25044 32212
rect 25038 32172 25044 32184
rect 25096 32172 25102 32224
rect 26206 32212 26234 32252
rect 27982 32240 27988 32292
rect 28040 32280 28046 32292
rect 28629 32283 28687 32289
rect 28629 32280 28641 32283
rect 28040 32252 28641 32280
rect 28040 32240 28046 32252
rect 28629 32249 28641 32252
rect 28675 32280 28687 32283
rect 28718 32280 28724 32292
rect 28675 32252 28724 32280
rect 28675 32249 28687 32252
rect 28629 32243 28687 32249
rect 28718 32240 28724 32252
rect 28776 32240 28782 32292
rect 31110 32212 31116 32224
rect 26206 32184 31116 32212
rect 31110 32172 31116 32184
rect 31168 32172 31174 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 10410 32008 10416 32020
rect 10371 31980 10416 32008
rect 10410 31968 10416 31980
rect 10468 31968 10474 32020
rect 12158 31968 12164 32020
rect 12216 32008 12222 32020
rect 19610 32008 19616 32020
rect 12216 31980 13584 32008
rect 19571 31980 19616 32008
rect 12216 31968 12222 31980
rect 4433 31943 4491 31949
rect 4433 31909 4445 31943
rect 4479 31940 4491 31943
rect 4798 31940 4804 31952
rect 4479 31912 4804 31940
rect 4479 31909 4491 31912
rect 4433 31903 4491 31909
rect 4798 31900 4804 31912
rect 4856 31900 4862 31952
rect 8938 31832 8944 31884
rect 8996 31872 9002 31884
rect 10229 31875 10287 31881
rect 8996 31844 10180 31872
rect 8996 31832 9002 31844
rect 1578 31764 1584 31816
rect 1636 31804 1642 31816
rect 1673 31807 1731 31813
rect 1673 31804 1685 31807
rect 1636 31776 1685 31804
rect 1636 31764 1642 31776
rect 1673 31773 1685 31776
rect 1719 31773 1731 31807
rect 2498 31804 2504 31816
rect 2459 31776 2504 31804
rect 1673 31767 1731 31773
rect 2498 31764 2504 31776
rect 2556 31764 2562 31816
rect 4617 31807 4675 31813
rect 4617 31773 4629 31807
rect 4663 31804 4675 31807
rect 9950 31804 9956 31816
rect 4663 31776 9956 31804
rect 4663 31773 4675 31776
rect 4617 31767 4675 31773
rect 9950 31764 9956 31776
rect 10008 31764 10014 31816
rect 10152 31813 10180 31844
rect 10229 31841 10241 31875
rect 10275 31872 10287 31875
rect 11790 31872 11796 31884
rect 10275 31844 11796 31872
rect 10275 31841 10287 31844
rect 10229 31835 10287 31841
rect 11790 31832 11796 31844
rect 11848 31832 11854 31884
rect 13556 31881 13584 31980
rect 19610 31968 19616 31980
rect 19668 31968 19674 32020
rect 19794 31968 19800 32020
rect 19852 32008 19858 32020
rect 20622 32008 20628 32020
rect 19852 31980 20628 32008
rect 19852 31968 19858 31980
rect 20622 31968 20628 31980
rect 20680 31968 20686 32020
rect 24765 32011 24823 32017
rect 24765 31977 24777 32011
rect 24811 32008 24823 32011
rect 24854 32008 24860 32020
rect 24811 31980 24860 32008
rect 24811 31977 24823 31980
rect 24765 31971 24823 31977
rect 24854 31968 24860 31980
rect 24912 31968 24918 32020
rect 24949 32011 25007 32017
rect 24949 31977 24961 32011
rect 24995 32008 25007 32011
rect 25314 32008 25320 32020
rect 24995 31980 25320 32008
rect 24995 31977 25007 31980
rect 24949 31971 25007 31977
rect 25314 31968 25320 31980
rect 25372 31968 25378 32020
rect 27062 32008 27068 32020
rect 27023 31980 27068 32008
rect 27062 31968 27068 31980
rect 27120 31968 27126 32020
rect 27893 32011 27951 32017
rect 27893 31977 27905 32011
rect 27939 32008 27951 32011
rect 27982 32008 27988 32020
rect 27939 31980 27988 32008
rect 27939 31977 27951 31980
rect 27893 31971 27951 31977
rect 27982 31968 27988 31980
rect 28040 31968 28046 32020
rect 28534 32008 28540 32020
rect 28495 31980 28540 32008
rect 28534 31968 28540 31980
rect 28592 31968 28598 32020
rect 31110 32008 31116 32020
rect 31071 31980 31116 32008
rect 31110 31968 31116 31980
rect 31168 31968 31174 32020
rect 13906 31900 13912 31952
rect 13964 31940 13970 31952
rect 14918 31940 14924 31952
rect 13964 31912 14924 31940
rect 13964 31900 13970 31912
rect 14918 31900 14924 31912
rect 14976 31940 14982 31952
rect 15013 31943 15071 31949
rect 15013 31940 15025 31943
rect 14976 31912 15025 31940
rect 14976 31900 14982 31912
rect 15013 31909 15025 31912
rect 15059 31940 15071 31943
rect 18141 31943 18199 31949
rect 15059 31912 17080 31940
rect 15059 31909 15071 31912
rect 15013 31903 15071 31909
rect 13541 31875 13599 31881
rect 13541 31841 13553 31875
rect 13587 31872 13599 31875
rect 15194 31872 15200 31884
rect 13587 31844 15200 31872
rect 13587 31841 13599 31844
rect 13541 31835 13599 31841
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 16022 31832 16028 31884
rect 16080 31872 16086 31884
rect 16945 31875 17003 31881
rect 16945 31872 16957 31875
rect 16080 31844 16957 31872
rect 16080 31832 16086 31844
rect 16945 31841 16957 31844
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 10137 31807 10195 31813
rect 10137 31773 10149 31807
rect 10183 31773 10195 31807
rect 13285 31807 13343 31813
rect 10137 31767 10195 31773
rect 10244 31776 12204 31804
rect 9398 31736 9404 31748
rect 9311 31708 9404 31736
rect 9398 31696 9404 31708
rect 9456 31736 9462 31748
rect 10244 31736 10272 31776
rect 9456 31708 10272 31736
rect 9456 31696 9462 31708
rect 1762 31628 1768 31680
rect 1820 31668 1826 31680
rect 2409 31671 2467 31677
rect 2409 31668 2421 31671
rect 1820 31640 2421 31668
rect 1820 31628 1826 31640
rect 2409 31637 2421 31640
rect 2455 31637 2467 31671
rect 9306 31668 9312 31680
rect 9267 31640 9312 31668
rect 2409 31631 2467 31637
rect 9306 31628 9312 31640
rect 9364 31628 9370 31680
rect 12176 31677 12204 31776
rect 13285 31773 13297 31807
rect 13331 31804 13343 31807
rect 14274 31804 14280 31816
rect 13331 31776 14280 31804
rect 13331 31773 13343 31776
rect 13285 31767 13343 31773
rect 14274 31764 14280 31776
rect 14332 31764 14338 31816
rect 15381 31807 15439 31813
rect 15381 31804 15393 31807
rect 14384 31776 15393 31804
rect 13538 31696 13544 31748
rect 13596 31736 13602 31748
rect 14384 31736 14412 31776
rect 15381 31773 15393 31776
rect 15427 31773 15439 31807
rect 15381 31767 15439 31773
rect 15565 31807 15623 31813
rect 15565 31773 15577 31807
rect 15611 31804 15623 31807
rect 16666 31804 16672 31816
rect 15611 31776 16672 31804
rect 15611 31773 15623 31776
rect 15565 31767 15623 31773
rect 16666 31764 16672 31776
rect 16724 31764 16730 31816
rect 16761 31807 16819 31813
rect 16761 31773 16773 31807
rect 16807 31804 16819 31807
rect 17052 31804 17080 31912
rect 18141 31909 18153 31943
rect 18187 31940 18199 31943
rect 18187 31912 21128 31940
rect 18187 31909 18199 31912
rect 18141 31903 18199 31909
rect 20254 31872 20260 31884
rect 19536 31844 20260 31872
rect 17586 31804 17592 31816
rect 16807 31776 17592 31804
rect 16807 31773 16819 31776
rect 16761 31767 16819 31773
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 18322 31764 18328 31816
rect 18380 31804 18386 31816
rect 19536 31813 19564 31844
rect 20254 31832 20260 31844
rect 20312 31832 20318 31884
rect 20530 31872 20536 31884
rect 20491 31844 20536 31872
rect 20530 31832 20536 31844
rect 20588 31832 20594 31884
rect 20622 31832 20628 31884
rect 20680 31872 20686 31884
rect 20901 31875 20959 31881
rect 20680 31844 20725 31872
rect 20680 31832 20686 31844
rect 20901 31841 20913 31875
rect 20947 31872 20959 31875
rect 20990 31872 20996 31884
rect 20947 31844 20996 31872
rect 20947 31841 20959 31844
rect 20901 31835 20959 31841
rect 20990 31832 20996 31844
rect 21048 31832 21054 31884
rect 18417 31807 18475 31813
rect 18417 31804 18429 31807
rect 18380 31776 18429 31804
rect 18380 31764 18386 31776
rect 18417 31773 18429 31776
rect 18463 31773 18475 31807
rect 19521 31807 19579 31813
rect 19521 31804 19533 31807
rect 18417 31767 18475 31773
rect 19260 31776 19533 31804
rect 15289 31739 15347 31745
rect 15289 31736 15301 31739
rect 13596 31708 14412 31736
rect 15028 31708 15301 31736
rect 13596 31696 13602 31708
rect 12161 31671 12219 31677
rect 12161 31637 12173 31671
rect 12207 31668 12219 31671
rect 15028 31668 15056 31708
rect 15289 31705 15301 31708
rect 15335 31705 15347 31739
rect 18138 31736 18144 31748
rect 18099 31708 18144 31736
rect 15289 31699 15347 31705
rect 18138 31696 18144 31708
rect 18196 31696 18202 31748
rect 12207 31640 15056 31668
rect 15197 31671 15255 31677
rect 12207 31637 12219 31640
rect 12161 31631 12219 31637
rect 15197 31637 15209 31671
rect 15243 31668 15255 31671
rect 15378 31668 15384 31680
rect 15243 31640 15384 31668
rect 15243 31637 15255 31640
rect 15197 31631 15255 31637
rect 15378 31628 15384 31640
rect 15436 31668 15442 31680
rect 15654 31668 15660 31680
rect 15436 31640 15660 31668
rect 15436 31628 15442 31640
rect 15654 31628 15660 31640
rect 15712 31628 15718 31680
rect 18325 31671 18383 31677
rect 18325 31637 18337 31671
rect 18371 31668 18383 31671
rect 18414 31668 18420 31680
rect 18371 31640 18420 31668
rect 18371 31637 18383 31640
rect 18325 31631 18383 31637
rect 18414 31628 18420 31640
rect 18472 31668 18478 31680
rect 19260 31668 19288 31776
rect 19521 31773 19533 31776
rect 19567 31773 19579 31807
rect 19521 31767 19579 31773
rect 19705 31807 19763 31813
rect 19705 31773 19717 31807
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 19720 31736 19748 31767
rect 19794 31764 19800 31816
rect 19852 31804 19858 31816
rect 20441 31807 20499 31813
rect 20441 31804 20453 31807
rect 19852 31776 19897 31804
rect 20364 31776 20453 31804
rect 19852 31764 19858 31776
rect 20070 31736 20076 31748
rect 19720 31708 20076 31736
rect 20070 31696 20076 31708
rect 20128 31696 20134 31748
rect 18472 31640 19288 31668
rect 18472 31628 18478 31640
rect 19334 31628 19340 31680
rect 19392 31668 19398 31680
rect 20364 31668 20392 31776
rect 20441 31773 20453 31776
rect 20487 31773 20499 31807
rect 20441 31767 20499 31773
rect 20717 31807 20775 31813
rect 20717 31773 20729 31807
rect 20763 31804 20775 31807
rect 20806 31804 20812 31816
rect 20763 31776 20812 31804
rect 20763 31773 20775 31776
rect 20717 31767 20775 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 21100 31804 21128 31912
rect 22462 31900 22468 31952
rect 22520 31940 22526 31952
rect 22833 31943 22891 31949
rect 22833 31940 22845 31943
rect 22520 31912 22845 31940
rect 22520 31900 22526 31912
rect 22833 31909 22845 31912
rect 22879 31940 22891 31943
rect 22879 31912 23704 31940
rect 22879 31909 22891 31912
rect 22833 31903 22891 31909
rect 21450 31872 21456 31884
rect 21411 31844 21456 31872
rect 21450 31832 21456 31844
rect 21508 31832 21514 31884
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31841 23627 31875
rect 23676 31872 23704 31912
rect 25222 31900 25228 31952
rect 25280 31940 25286 31952
rect 27709 31943 27767 31949
rect 27709 31940 27721 31943
rect 25280 31912 27721 31940
rect 25280 31900 25286 31912
rect 27709 31909 27721 31912
rect 27755 31909 27767 31943
rect 27709 31903 27767 31909
rect 26970 31872 26976 31884
rect 23676 31844 26976 31872
rect 23569 31835 23627 31841
rect 21709 31807 21767 31813
rect 21709 31804 21721 31807
rect 21100 31776 21721 31804
rect 21709 31773 21721 31776
rect 21755 31773 21767 31807
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 21709 31767 21767 31773
rect 21836 31776 23489 31804
rect 20530 31696 20536 31748
rect 20588 31736 20594 31748
rect 21836 31736 21864 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23584 31804 23612 31835
rect 26970 31832 26976 31844
rect 27028 31832 27034 31884
rect 27157 31875 27215 31881
rect 27157 31841 27169 31875
rect 27203 31872 27215 31875
rect 27798 31872 27804 31884
rect 27203 31844 27804 31872
rect 27203 31841 27215 31844
rect 27157 31835 27215 31841
rect 27798 31832 27804 31844
rect 27856 31872 27862 31884
rect 27856 31844 28580 31872
rect 27856 31832 27862 31844
rect 25498 31804 25504 31816
rect 23584 31776 25504 31804
rect 23477 31767 23535 31773
rect 25498 31764 25504 31776
rect 25556 31764 25562 31816
rect 27249 31807 27307 31813
rect 27249 31773 27261 31807
rect 27295 31804 27307 31807
rect 28258 31804 28264 31816
rect 27295 31776 28264 31804
rect 27295 31773 27307 31776
rect 27249 31767 27307 31773
rect 28258 31764 28264 31776
rect 28316 31764 28322 31816
rect 28552 31813 28580 31844
rect 28537 31807 28595 31813
rect 28537 31773 28549 31807
rect 28583 31773 28595 31807
rect 28718 31804 28724 31816
rect 28679 31776 28724 31804
rect 28537 31767 28595 31773
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 29730 31804 29736 31816
rect 29691 31776 29736 31804
rect 29730 31764 29736 31776
rect 29788 31764 29794 31816
rect 33778 31804 33784 31816
rect 33739 31776 33784 31804
rect 33778 31764 33784 31776
rect 33836 31764 33842 31816
rect 20588 31708 21864 31736
rect 24581 31739 24639 31745
rect 20588 31696 20594 31708
rect 24581 31705 24593 31739
rect 24627 31705 24639 31739
rect 24581 31699 24639 31705
rect 19392 31640 20392 31668
rect 23845 31671 23903 31677
rect 19392 31628 19398 31640
rect 23845 31637 23857 31671
rect 23891 31668 23903 31671
rect 24394 31668 24400 31680
rect 23891 31640 24400 31668
rect 23891 31637 23903 31640
rect 23845 31631 23903 31637
rect 24394 31628 24400 31640
rect 24452 31668 24458 31680
rect 24596 31668 24624 31699
rect 27522 31696 27528 31748
rect 27580 31736 27586 31748
rect 27861 31739 27919 31745
rect 27861 31736 27873 31739
rect 27580 31708 27873 31736
rect 27580 31696 27586 31708
rect 27861 31705 27873 31708
rect 27907 31705 27919 31739
rect 28074 31736 28080 31748
rect 28035 31708 28080 31736
rect 27861 31699 27919 31705
rect 28074 31696 28080 31708
rect 28132 31696 28138 31748
rect 30000 31739 30058 31745
rect 30000 31705 30012 31739
rect 30046 31736 30058 31739
rect 30098 31736 30104 31748
rect 30046 31708 30104 31736
rect 30046 31705 30058 31708
rect 30000 31699 30058 31705
rect 30098 31696 30104 31708
rect 30156 31696 30162 31748
rect 24452 31640 24624 31668
rect 24452 31628 24458 31640
rect 24762 31628 24768 31680
rect 24820 31677 24826 31680
rect 24820 31671 24839 31677
rect 24827 31637 24839 31671
rect 24820 31631 24839 31637
rect 33873 31671 33931 31677
rect 33873 31637 33885 31671
rect 33919 31668 33931 31671
rect 34054 31668 34060 31680
rect 33919 31640 34060 31668
rect 33919 31637 33931 31640
rect 33873 31631 33931 31637
rect 24820 31628 24826 31631
rect 34054 31628 34060 31640
rect 34112 31628 34118 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 3513 31467 3571 31473
rect 3513 31433 3525 31467
rect 3559 31464 3571 31467
rect 3694 31464 3700 31476
rect 3559 31436 3700 31464
rect 3559 31433 3571 31436
rect 3513 31427 3571 31433
rect 3694 31424 3700 31436
rect 3752 31424 3758 31476
rect 6886 31436 12434 31464
rect 6886 31396 6914 31436
rect 2332 31368 6914 31396
rect 12406 31396 12434 31436
rect 14182 31424 14188 31476
rect 14240 31464 14246 31476
rect 14645 31467 14703 31473
rect 14645 31464 14657 31467
rect 14240 31436 14657 31464
rect 14240 31424 14246 31436
rect 14645 31433 14657 31436
rect 14691 31433 14703 31467
rect 18138 31464 18144 31476
rect 14645 31427 14703 31433
rect 14752 31436 16620 31464
rect 18099 31436 18144 31464
rect 14752 31396 14780 31436
rect 12406 31368 14780 31396
rect 14829 31399 14887 31405
rect 2332 31340 2360 31368
rect 14829 31365 14841 31399
rect 14875 31396 14887 31399
rect 15657 31399 15715 31405
rect 15657 31396 15669 31399
rect 14875 31368 15669 31396
rect 14875 31365 14887 31368
rect 14829 31359 14887 31365
rect 15657 31365 15669 31368
rect 15703 31365 15715 31399
rect 16592 31396 16620 31436
rect 18138 31424 18144 31436
rect 18196 31424 18202 31476
rect 24581 31467 24639 31473
rect 24581 31433 24593 31467
rect 24627 31464 24639 31467
rect 24946 31464 24952 31476
rect 24627 31436 24952 31464
rect 24627 31433 24639 31436
rect 24581 31427 24639 31433
rect 24946 31424 24952 31436
rect 25004 31424 25010 31476
rect 25130 31464 25136 31476
rect 25091 31436 25136 31464
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 26234 31464 26240 31476
rect 26195 31436 26240 31464
rect 26234 31424 26240 31436
rect 26292 31424 26298 31476
rect 27801 31467 27859 31473
rect 27801 31433 27813 31467
rect 27847 31464 27859 31467
rect 28074 31464 28080 31476
rect 27847 31436 28080 31464
rect 27847 31433 27859 31436
rect 27801 31427 27859 31433
rect 28074 31424 28080 31436
rect 28132 31424 28138 31476
rect 30098 31464 30104 31476
rect 30059 31436 30104 31464
rect 30098 31424 30104 31436
rect 30156 31424 30162 31476
rect 20714 31396 20720 31408
rect 15657 31359 15715 31365
rect 15764 31368 16160 31396
rect 16592 31368 20720 31396
rect 2314 31328 2320 31340
rect 2275 31300 2320 31328
rect 2314 31288 2320 31300
rect 2372 31288 2378 31340
rect 3602 31328 3608 31340
rect 3563 31300 3608 31328
rect 3602 31288 3608 31300
rect 3660 31288 3666 31340
rect 9030 31288 9036 31340
rect 9088 31328 9094 31340
rect 9493 31331 9551 31337
rect 9493 31328 9505 31331
rect 9088 31300 9505 31328
rect 9088 31288 9094 31300
rect 9493 31297 9505 31300
rect 9539 31297 9551 31331
rect 9674 31328 9680 31340
rect 9635 31300 9680 31328
rect 9493 31291 9551 31297
rect 9674 31288 9680 31300
rect 9732 31288 9738 31340
rect 15102 31288 15108 31340
rect 15160 31328 15166 31340
rect 15764 31328 15792 31368
rect 15160 31300 15792 31328
rect 15160 31288 15166 31300
rect 15838 31288 15844 31340
rect 15896 31328 15902 31340
rect 16022 31328 16028 31340
rect 15896 31300 15941 31328
rect 15983 31300 16028 31328
rect 15896 31288 15902 31300
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 16132 31337 16160 31368
rect 20714 31356 20720 31368
rect 20772 31356 20778 31408
rect 24854 31356 24860 31408
rect 24912 31396 24918 31408
rect 25961 31399 26019 31405
rect 25961 31396 25973 31399
rect 24912 31368 25973 31396
rect 24912 31356 24918 31368
rect 25961 31365 25973 31368
rect 26007 31396 26019 31399
rect 26142 31396 26148 31408
rect 26007 31368 26148 31396
rect 26007 31365 26019 31368
rect 25961 31359 26019 31365
rect 26142 31356 26148 31368
rect 26200 31356 26206 31408
rect 27246 31396 27252 31408
rect 26252 31368 27252 31396
rect 26252 31340 26280 31368
rect 27246 31356 27252 31368
rect 27304 31356 27310 31408
rect 34054 31396 34060 31408
rect 34015 31368 34060 31396
rect 34054 31356 34060 31368
rect 34112 31356 34118 31408
rect 35710 31396 35716 31408
rect 35671 31368 35716 31396
rect 35710 31356 35716 31368
rect 35768 31356 35774 31408
rect 16117 31331 16175 31337
rect 16117 31297 16129 31331
rect 16163 31297 16175 31331
rect 18414 31328 18420 31340
rect 18375 31300 18420 31328
rect 16117 31291 16175 31297
rect 18414 31288 18420 31300
rect 18472 31288 18478 31340
rect 24394 31328 24400 31340
rect 24355 31300 24400 31328
rect 24394 31288 24400 31300
rect 24452 31288 24458 31340
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31328 24639 31331
rect 24670 31328 24676 31340
rect 24627 31300 24676 31328
rect 24627 31297 24639 31300
rect 24581 31291 24639 31297
rect 8570 31260 8576 31272
rect 8483 31232 8576 31260
rect 8570 31220 8576 31232
rect 8628 31260 8634 31272
rect 9306 31260 9312 31272
rect 8628 31232 9312 31260
rect 8628 31220 8634 31232
rect 9306 31220 9312 31232
rect 9364 31220 9370 31272
rect 11054 31220 11060 31272
rect 11112 31260 11118 31272
rect 11698 31260 11704 31272
rect 11112 31232 11704 31260
rect 11112 31220 11118 31232
rect 11698 31220 11704 31232
rect 11756 31260 11762 31272
rect 17218 31260 17224 31272
rect 11756 31232 17224 31260
rect 11756 31220 11762 31232
rect 17218 31220 17224 31232
rect 17276 31220 17282 31272
rect 18046 31220 18052 31272
rect 18104 31260 18110 31272
rect 18141 31263 18199 31269
rect 18141 31260 18153 31263
rect 18104 31232 18153 31260
rect 18104 31220 18110 31232
rect 18141 31229 18153 31232
rect 18187 31229 18199 31263
rect 18322 31260 18328 31272
rect 18283 31232 18328 31260
rect 18141 31223 18199 31229
rect 18322 31220 18328 31232
rect 18380 31220 18386 31272
rect 21174 31220 21180 31272
rect 21232 31260 21238 31272
rect 24596 31260 24624 31291
rect 24670 31288 24676 31300
rect 24728 31288 24734 31340
rect 25038 31328 25044 31340
rect 24999 31300 25044 31328
rect 25038 31288 25044 31300
rect 25096 31288 25102 31340
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31328 25283 31331
rect 25590 31328 25596 31340
rect 25271 31300 25596 31328
rect 25271 31297 25283 31300
rect 25225 31291 25283 31297
rect 25590 31288 25596 31300
rect 25648 31288 25654 31340
rect 25866 31328 25872 31340
rect 25827 31300 25872 31328
rect 25866 31288 25872 31300
rect 25924 31288 25930 31340
rect 26053 31331 26111 31337
rect 26053 31297 26065 31331
rect 26099 31328 26111 31331
rect 26234 31328 26240 31340
rect 26099 31300 26240 31328
rect 26099 31297 26111 31300
rect 26053 31291 26111 31297
rect 26234 31288 26240 31300
rect 26292 31288 26298 31340
rect 26970 31288 26976 31340
rect 27028 31328 27034 31340
rect 27433 31331 27491 31337
rect 27433 31328 27445 31331
rect 27028 31300 27445 31328
rect 27028 31288 27034 31300
rect 27433 31297 27445 31300
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 30009 31331 30067 31337
rect 30009 31297 30021 31331
rect 30055 31297 30067 31331
rect 30009 31291 30067 31297
rect 30193 31331 30251 31337
rect 30193 31297 30205 31331
rect 30239 31328 30251 31331
rect 30558 31328 30564 31340
rect 30239 31300 30564 31328
rect 30239 31297 30251 31300
rect 30193 31291 30251 31297
rect 21232 31232 24624 31260
rect 27525 31263 27583 31269
rect 21232 31220 21238 31232
rect 27525 31229 27537 31263
rect 27571 31260 27583 31263
rect 28166 31260 28172 31272
rect 27571 31232 28172 31260
rect 27571 31229 27583 31232
rect 27525 31223 27583 31229
rect 28166 31220 28172 31232
rect 28224 31260 28230 31272
rect 28902 31260 28908 31272
rect 28224 31232 28908 31260
rect 28224 31220 28230 31232
rect 28902 31220 28908 31232
rect 28960 31220 28966 31272
rect 30024 31260 30052 31291
rect 30558 31288 30564 31300
rect 30616 31288 30622 31340
rect 33870 31260 33876 31272
rect 30024 31232 33876 31260
rect 33870 31220 33876 31232
rect 33928 31220 33934 31272
rect 2225 31195 2283 31201
rect 2225 31161 2237 31195
rect 2271 31192 2283 31195
rect 3234 31192 3240 31204
rect 2271 31164 3240 31192
rect 2271 31161 2283 31164
rect 2225 31155 2283 31161
rect 3234 31152 3240 31164
rect 3292 31152 3298 31204
rect 8938 31192 8944 31204
rect 8899 31164 8944 31192
rect 8938 31152 8944 31164
rect 8996 31152 9002 31204
rect 15197 31195 15255 31201
rect 15197 31161 15209 31195
rect 15243 31192 15255 31195
rect 15286 31192 15292 31204
rect 15243 31164 15292 31192
rect 15243 31161 15255 31164
rect 15197 31155 15255 31161
rect 15286 31152 15292 31164
rect 15344 31152 15350 31204
rect 25685 31195 25743 31201
rect 25685 31161 25697 31195
rect 25731 31192 25743 31195
rect 26694 31192 26700 31204
rect 25731 31164 26700 31192
rect 25731 31161 25743 31164
rect 25685 31155 25743 31161
rect 26694 31152 26700 31164
rect 26752 31192 26758 31204
rect 27338 31192 27344 31204
rect 26752 31164 27344 31192
rect 26752 31152 26758 31164
rect 27338 31152 27344 31164
rect 27396 31152 27402 31204
rect 2958 31124 2964 31136
rect 2919 31096 2964 31124
rect 2958 31084 2964 31096
rect 3016 31084 3022 31136
rect 4062 31124 4068 31136
rect 4023 31096 4068 31124
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 9030 31124 9036 31136
rect 8991 31096 9036 31124
rect 9030 31084 9036 31096
rect 9088 31084 9094 31136
rect 9490 31124 9496 31136
rect 9451 31096 9496 31124
rect 9490 31084 9496 31096
rect 9548 31084 9554 31136
rect 14734 31084 14740 31136
rect 14792 31124 14798 31136
rect 14829 31127 14887 31133
rect 14829 31124 14841 31127
rect 14792 31096 14841 31124
rect 14792 31084 14798 31096
rect 14829 31093 14841 31096
rect 14875 31093 14887 31127
rect 14829 31087 14887 31093
rect 15010 31084 15016 31136
rect 15068 31124 15074 31136
rect 19426 31124 19432 31136
rect 15068 31096 19432 31124
rect 15068 31084 15074 31096
rect 19426 31084 19432 31096
rect 19484 31124 19490 31136
rect 20530 31124 20536 31136
rect 19484 31096 20536 31124
rect 19484 31084 19490 31096
rect 20530 31084 20536 31096
rect 20588 31084 20594 31136
rect 37829 31127 37887 31133
rect 37829 31093 37841 31127
rect 37875 31124 37887 31127
rect 38286 31124 38292 31136
rect 37875 31096 38292 31124
rect 37875 31093 37887 31096
rect 37829 31087 37887 31093
rect 38286 31084 38292 31096
rect 38344 31084 38350 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 3602 30880 3608 30932
rect 3660 30920 3666 30932
rect 4525 30923 4583 30929
rect 4525 30920 4537 30923
rect 3660 30892 4537 30920
rect 3660 30880 3666 30892
rect 4525 30889 4537 30892
rect 4571 30889 4583 30923
rect 14274 30920 14280 30932
rect 14235 30892 14280 30920
rect 4525 30883 4583 30889
rect 14274 30880 14280 30892
rect 14332 30880 14338 30932
rect 15838 30920 15844 30932
rect 14568 30892 15844 30920
rect 13541 30855 13599 30861
rect 13541 30821 13553 30855
rect 13587 30852 13599 30855
rect 14568 30852 14596 30892
rect 15838 30880 15844 30892
rect 15896 30880 15902 30932
rect 17218 30880 17224 30932
rect 17276 30920 17282 30932
rect 22373 30923 22431 30929
rect 17276 30892 22094 30920
rect 17276 30880 17282 30892
rect 13587 30824 14596 30852
rect 14645 30855 14703 30861
rect 13587 30821 13599 30824
rect 13541 30815 13599 30821
rect 14645 30821 14657 30855
rect 14691 30852 14703 30855
rect 15286 30852 15292 30864
rect 14691 30824 15292 30852
rect 14691 30821 14703 30824
rect 14645 30815 14703 30821
rect 15286 30812 15292 30824
rect 15344 30812 15350 30864
rect 20622 30852 20628 30864
rect 17236 30824 20628 30852
rect 1578 30784 1584 30796
rect 1539 30756 1584 30784
rect 1578 30744 1584 30756
rect 1636 30744 1642 30796
rect 1762 30784 1768 30796
rect 1723 30756 1768 30784
rect 1762 30744 1768 30756
rect 1820 30744 1826 30796
rect 2774 30784 2780 30796
rect 2735 30756 2780 30784
rect 2774 30744 2780 30756
rect 2832 30744 2838 30796
rect 9306 30744 9312 30796
rect 9364 30784 9370 30796
rect 13725 30787 13783 30793
rect 9364 30756 13676 30784
rect 9364 30744 9370 30756
rect 10134 30676 10140 30728
rect 10192 30716 10198 30728
rect 10781 30719 10839 30725
rect 10781 30716 10793 30719
rect 10192 30688 10793 30716
rect 10192 30676 10198 30688
rect 10781 30685 10793 30688
rect 10827 30685 10839 30719
rect 11054 30716 11060 30728
rect 11015 30688 11060 30716
rect 10781 30679 10839 30685
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 13354 30676 13360 30728
rect 13412 30716 13418 30728
rect 13449 30719 13507 30725
rect 13449 30716 13461 30719
rect 13412 30688 13461 30716
rect 13412 30676 13418 30688
rect 13449 30685 13461 30688
rect 13495 30685 13507 30719
rect 13648 30716 13676 30756
rect 13725 30753 13737 30787
rect 13771 30784 13783 30787
rect 14274 30784 14280 30796
rect 13771 30756 14280 30784
rect 13771 30753 13783 30756
rect 13725 30747 13783 30753
rect 14274 30744 14280 30756
rect 14332 30744 14338 30796
rect 14737 30787 14795 30793
rect 14737 30784 14749 30787
rect 14384 30756 14749 30784
rect 14384 30716 14412 30756
rect 14737 30753 14749 30756
rect 14783 30784 14795 30787
rect 15010 30784 15016 30796
rect 14783 30756 15016 30784
rect 14783 30753 14795 30756
rect 14737 30747 14795 30753
rect 15010 30744 15016 30756
rect 15068 30744 15074 30796
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 15657 30787 15715 30793
rect 15657 30784 15669 30787
rect 15252 30756 15669 30784
rect 15252 30744 15258 30756
rect 15657 30753 15669 30756
rect 15703 30753 15715 30787
rect 15657 30747 15715 30753
rect 13648 30688 14412 30716
rect 14461 30719 14519 30725
rect 13449 30679 13507 30685
rect 14461 30685 14473 30719
rect 14507 30685 14519 30719
rect 14461 30679 14519 30685
rect 4433 30651 4491 30657
rect 4433 30617 4445 30651
rect 4479 30617 4491 30651
rect 14476 30648 14504 30679
rect 17236 30648 17264 30824
rect 20622 30812 20628 30824
rect 20680 30812 20686 30864
rect 22066 30852 22094 30892
rect 22373 30889 22385 30923
rect 22419 30920 22431 30923
rect 25038 30920 25044 30932
rect 22419 30892 25044 30920
rect 22419 30889 22431 30892
rect 22373 30883 22431 30889
rect 25038 30880 25044 30892
rect 25096 30880 25102 30932
rect 25590 30920 25596 30932
rect 25551 30892 25596 30920
rect 25590 30880 25596 30892
rect 25648 30880 25654 30932
rect 26510 30920 26516 30932
rect 25700 30892 26516 30920
rect 25700 30852 25728 30892
rect 26510 30880 26516 30892
rect 26568 30880 26574 30932
rect 27801 30923 27859 30929
rect 27801 30889 27813 30923
rect 27847 30920 27859 30923
rect 28258 30920 28264 30932
rect 27847 30892 28264 30920
rect 27847 30889 27859 30892
rect 27801 30883 27859 30889
rect 28258 30880 28264 30892
rect 28316 30880 28322 30932
rect 28902 30880 28908 30932
rect 28960 30920 28966 30932
rect 30101 30923 30159 30929
rect 30101 30920 30113 30923
rect 28960 30892 30113 30920
rect 28960 30880 28966 30892
rect 30101 30889 30113 30892
rect 30147 30889 30159 30923
rect 30101 30883 30159 30889
rect 26694 30852 26700 30864
rect 22066 30824 25728 30852
rect 25884 30824 26700 30852
rect 25884 30796 25912 30824
rect 26694 30812 26700 30824
rect 26752 30812 26758 30864
rect 18690 30784 18696 30796
rect 17972 30756 18696 30784
rect 17972 30728 18000 30756
rect 18690 30744 18696 30756
rect 18748 30744 18754 30796
rect 19058 30744 19064 30796
rect 19116 30784 19122 30796
rect 19429 30787 19487 30793
rect 19429 30784 19441 30787
rect 19116 30756 19441 30784
rect 19116 30744 19122 30756
rect 19429 30753 19441 30756
rect 19475 30753 19487 30787
rect 19429 30747 19487 30753
rect 19613 30787 19671 30793
rect 19613 30753 19625 30787
rect 19659 30784 19671 30787
rect 20438 30784 20444 30796
rect 19659 30756 20444 30784
rect 19659 30753 19671 30756
rect 19613 30747 19671 30753
rect 17310 30676 17316 30728
rect 17368 30716 17374 30728
rect 17865 30719 17923 30725
rect 17865 30716 17877 30719
rect 17368 30688 17877 30716
rect 17368 30676 17374 30688
rect 17865 30685 17877 30688
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 17954 30676 17960 30728
rect 18012 30716 18018 30728
rect 18141 30719 18199 30725
rect 18012 30688 18105 30716
rect 18012 30676 18018 30688
rect 18141 30685 18153 30719
rect 18187 30716 18199 30719
rect 18322 30716 18328 30728
rect 18187 30688 18328 30716
rect 18187 30685 18199 30688
rect 18141 30679 18199 30685
rect 18322 30676 18328 30688
rect 18380 30716 18386 30728
rect 18601 30719 18659 30725
rect 18601 30716 18613 30719
rect 18380 30688 18613 30716
rect 18380 30676 18386 30688
rect 18601 30685 18613 30688
rect 18647 30685 18659 30719
rect 18601 30679 18659 30685
rect 18785 30719 18843 30725
rect 18785 30685 18797 30719
rect 18831 30685 18843 30719
rect 18785 30679 18843 30685
rect 17402 30648 17408 30660
rect 14476 30620 17264 30648
rect 17363 30620 17408 30648
rect 4433 30611 4491 30617
rect 2866 30540 2872 30592
rect 2924 30580 2930 30592
rect 4448 30580 4476 30611
rect 17402 30608 17408 30620
rect 17460 30608 17466 30660
rect 18800 30648 18828 30679
rect 19334 30676 19340 30728
rect 19392 30716 19398 30728
rect 19628 30716 19656 30747
rect 20438 30744 20444 30756
rect 20496 30744 20502 30796
rect 25866 30784 25872 30796
rect 25827 30756 25872 30784
rect 25866 30744 25872 30756
rect 25924 30744 25930 30796
rect 26053 30787 26111 30793
rect 26053 30753 26065 30787
rect 26099 30784 26111 30787
rect 26142 30784 26148 30796
rect 26099 30756 26148 30784
rect 26099 30753 26111 30756
rect 26053 30747 26111 30753
rect 26142 30744 26148 30756
rect 26200 30744 26206 30796
rect 37826 30784 37832 30796
rect 37787 30756 37832 30784
rect 37826 30744 37832 30756
rect 37884 30744 37890 30796
rect 38286 30784 38292 30796
rect 38247 30756 38292 30784
rect 38286 30744 38292 30756
rect 38344 30744 38350 30796
rect 19392 30688 19656 30716
rect 19705 30719 19763 30725
rect 19392 30676 19398 30688
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 20070 30716 20076 30728
rect 19751 30688 20076 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 20070 30676 20076 30688
rect 20128 30676 20134 30728
rect 22094 30676 22100 30728
rect 22152 30716 22158 30728
rect 25777 30719 25835 30725
rect 22152 30688 22197 30716
rect 22152 30676 22158 30688
rect 25777 30685 25789 30719
rect 25823 30685 25835 30719
rect 25777 30679 25835 30685
rect 25961 30719 26019 30725
rect 25961 30685 25973 30719
rect 26007 30716 26019 30719
rect 26786 30716 26792 30728
rect 26007 30688 26792 30716
rect 26007 30685 26019 30688
rect 25961 30679 26019 30685
rect 19429 30651 19487 30657
rect 19429 30648 19441 30651
rect 18800 30620 19441 30648
rect 19429 30617 19441 30620
rect 19475 30617 19487 30651
rect 22370 30648 22376 30660
rect 22331 30620 22376 30648
rect 19429 30611 19487 30617
rect 22370 30608 22376 30620
rect 22428 30608 22434 30660
rect 25792 30648 25820 30679
rect 26786 30676 26792 30688
rect 26844 30716 26850 30728
rect 27246 30716 27252 30728
rect 26844 30688 27252 30716
rect 26844 30676 26850 30688
rect 27246 30676 27252 30688
rect 27304 30676 27310 30728
rect 27614 30716 27620 30728
rect 27575 30688 27620 30716
rect 27614 30676 27620 30688
rect 27672 30676 27678 30728
rect 27801 30719 27859 30725
rect 27801 30685 27813 30719
rect 27847 30685 27859 30719
rect 27801 30679 27859 30685
rect 26234 30648 26240 30660
rect 25792 30620 26240 30648
rect 26234 30608 26240 30620
rect 26292 30608 26298 30660
rect 27816 30648 27844 30679
rect 28626 30648 28632 30660
rect 27816 30620 28632 30648
rect 28626 30608 28632 30620
rect 28684 30648 28690 30660
rect 30009 30651 30067 30657
rect 30009 30648 30021 30651
rect 28684 30620 30021 30648
rect 28684 30608 28690 30620
rect 30009 30617 30021 30620
rect 30055 30617 30067 30651
rect 38102 30648 38108 30660
rect 38063 30620 38108 30648
rect 30009 30611 30067 30617
rect 38102 30608 38108 30620
rect 38160 30608 38166 30660
rect 13722 30580 13728 30592
rect 2924 30552 4476 30580
rect 13683 30552 13728 30580
rect 2924 30540 2930 30552
rect 13722 30540 13728 30552
rect 13780 30540 13786 30592
rect 18049 30583 18107 30589
rect 18049 30549 18061 30583
rect 18095 30580 18107 30583
rect 18230 30580 18236 30592
rect 18095 30552 18236 30580
rect 18095 30549 18107 30552
rect 18049 30543 18107 30549
rect 18230 30540 18236 30552
rect 18288 30540 18294 30592
rect 18690 30580 18696 30592
rect 18651 30552 18696 30580
rect 18690 30540 18696 30552
rect 18748 30540 18754 30592
rect 22189 30583 22247 30589
rect 22189 30549 22201 30583
rect 22235 30580 22247 30583
rect 23106 30580 23112 30592
rect 22235 30552 23112 30580
rect 22235 30549 22247 30552
rect 22189 30543 22247 30549
rect 23106 30540 23112 30552
rect 23164 30540 23170 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 15194 30376 15200 30388
rect 15155 30348 15200 30376
rect 15194 30336 15200 30348
rect 15252 30336 15258 30388
rect 15365 30379 15423 30385
rect 15365 30345 15377 30379
rect 15411 30376 15423 30379
rect 15838 30376 15844 30388
rect 15411 30348 15844 30376
rect 15411 30345 15423 30348
rect 15365 30339 15423 30345
rect 15838 30336 15844 30348
rect 15896 30336 15902 30388
rect 17310 30376 17316 30388
rect 17271 30348 17316 30376
rect 17310 30336 17316 30348
rect 17368 30336 17374 30388
rect 17402 30336 17408 30388
rect 17460 30376 17466 30388
rect 23382 30376 23388 30388
rect 17460 30348 23388 30376
rect 17460 30336 17466 30348
rect 23382 30336 23388 30348
rect 23440 30336 23446 30388
rect 26510 30336 26516 30388
rect 26568 30376 26574 30388
rect 27706 30376 27712 30388
rect 26568 30348 27712 30376
rect 26568 30336 26574 30348
rect 27706 30336 27712 30348
rect 27764 30336 27770 30388
rect 29730 30336 29736 30388
rect 29788 30336 29794 30388
rect 37645 30379 37703 30385
rect 37645 30345 37657 30379
rect 37691 30376 37703 30379
rect 38102 30376 38108 30388
rect 37691 30348 38108 30376
rect 37691 30345 37703 30348
rect 37645 30339 37703 30345
rect 38102 30336 38108 30348
rect 38160 30336 38166 30388
rect 9582 30308 9588 30320
rect 8772 30280 9588 30308
rect 2961 30243 3019 30249
rect 2961 30209 2973 30243
rect 3007 30240 3019 30243
rect 3142 30240 3148 30252
rect 3007 30212 3148 30240
rect 3007 30209 3019 30212
rect 2961 30203 3019 30209
rect 3142 30200 3148 30212
rect 3200 30200 3206 30252
rect 4062 30240 4068 30252
rect 4023 30212 4068 30240
rect 4062 30200 4068 30212
rect 4120 30200 4126 30252
rect 8113 30243 8171 30249
rect 8113 30209 8125 30243
rect 8159 30240 8171 30243
rect 8570 30240 8576 30252
rect 8159 30212 8576 30240
rect 8159 30209 8171 30212
rect 8113 30203 8171 30209
rect 8570 30200 8576 30212
rect 8628 30200 8634 30252
rect 8772 30249 8800 30280
rect 9582 30268 9588 30280
rect 9640 30308 9646 30320
rect 13722 30308 13728 30320
rect 9640 30280 13728 30308
rect 9640 30268 9646 30280
rect 13722 30268 13728 30280
rect 13780 30268 13786 30320
rect 15565 30311 15623 30317
rect 15565 30277 15577 30311
rect 15611 30308 15623 30311
rect 15654 30308 15660 30320
rect 15611 30280 15660 30308
rect 15611 30277 15623 30280
rect 15565 30271 15623 30277
rect 15654 30268 15660 30280
rect 15712 30308 15718 30320
rect 16022 30308 16028 30320
rect 15712 30280 16028 30308
rect 15712 30268 15718 30280
rect 16022 30268 16028 30280
rect 16080 30268 16086 30320
rect 16666 30268 16672 30320
rect 16724 30308 16730 30320
rect 17129 30311 17187 30317
rect 17129 30308 17141 30311
rect 16724 30280 17141 30308
rect 16724 30268 16730 30280
rect 17129 30277 17141 30280
rect 17175 30277 17187 30311
rect 17129 30271 17187 30277
rect 17221 30311 17279 30317
rect 17221 30277 17233 30311
rect 17267 30308 17279 30311
rect 17954 30308 17960 30320
rect 17267 30280 17960 30308
rect 17267 30277 17279 30280
rect 17221 30271 17279 30277
rect 8757 30243 8815 30249
rect 8757 30209 8769 30243
rect 8803 30209 8815 30243
rect 10134 30240 10140 30252
rect 10095 30212 10140 30240
rect 8757 30203 8815 30209
rect 10134 30200 10140 30212
rect 10192 30200 10198 30252
rect 11885 30243 11943 30249
rect 11885 30209 11897 30243
rect 11931 30240 11943 30243
rect 11974 30240 11980 30252
rect 11931 30212 11980 30240
rect 11931 30209 11943 30212
rect 11885 30203 11943 30209
rect 11974 30200 11980 30212
rect 12032 30200 12038 30252
rect 12069 30243 12127 30249
rect 12069 30209 12081 30243
rect 12115 30209 12127 30243
rect 12069 30203 12127 30209
rect 4249 30175 4307 30181
rect 4249 30141 4261 30175
rect 4295 30172 4307 30175
rect 4614 30172 4620 30184
rect 4295 30144 4620 30172
rect 4295 30141 4307 30144
rect 4249 30135 4307 30141
rect 4614 30132 4620 30144
rect 4672 30132 4678 30184
rect 4709 30175 4767 30181
rect 4709 30141 4721 30175
rect 4755 30141 4767 30175
rect 4709 30135 4767 30141
rect 8849 30175 8907 30181
rect 8849 30141 8861 30175
rect 8895 30172 8907 30175
rect 9490 30172 9496 30184
rect 8895 30144 9496 30172
rect 8895 30141 8907 30144
rect 8849 30135 8907 30141
rect 3050 30064 3056 30116
rect 3108 30104 3114 30116
rect 4724 30104 4752 30135
rect 9490 30132 9496 30144
rect 9548 30132 9554 30184
rect 9950 30132 9956 30184
rect 10008 30172 10014 30184
rect 10689 30175 10747 30181
rect 10689 30172 10701 30175
rect 10008 30144 10701 30172
rect 10008 30132 10014 30144
rect 10689 30141 10701 30144
rect 10735 30172 10747 30175
rect 12084 30172 12112 30203
rect 12158 30200 12164 30252
rect 12216 30240 12222 30252
rect 12216 30212 12261 30240
rect 12216 30200 12222 30212
rect 13078 30200 13084 30252
rect 13136 30240 13142 30252
rect 13538 30240 13544 30252
rect 13136 30212 13544 30240
rect 13136 30200 13142 30212
rect 13538 30200 13544 30212
rect 13596 30240 13602 30252
rect 14458 30240 14464 30252
rect 13596 30212 14464 30240
rect 13596 30200 13602 30212
rect 14458 30200 14464 30212
rect 14516 30240 14522 30252
rect 14553 30243 14611 30249
rect 14553 30240 14565 30243
rect 14516 30212 14565 30240
rect 14516 30200 14522 30212
rect 14553 30209 14565 30212
rect 14599 30209 14611 30243
rect 17144 30240 17172 30271
rect 17954 30268 17960 30280
rect 18012 30268 18018 30320
rect 18322 30308 18328 30320
rect 18283 30280 18328 30308
rect 18322 30268 18328 30280
rect 18380 30268 18386 30320
rect 19426 30308 19432 30320
rect 19387 30280 19432 30308
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 19521 30311 19579 30317
rect 19521 30277 19533 30311
rect 19567 30308 19579 30311
rect 19794 30308 19800 30320
rect 19567 30280 19800 30308
rect 19567 30277 19579 30280
rect 19521 30271 19579 30277
rect 19794 30268 19800 30280
rect 19852 30308 19858 30320
rect 23106 30308 23112 30320
rect 19852 30280 22094 30308
rect 23067 30280 23112 30308
rect 19852 30268 19858 30280
rect 18141 30243 18199 30249
rect 18141 30240 18153 30243
rect 17144 30212 18153 30240
rect 14553 30203 14611 30209
rect 18141 30209 18153 30212
rect 18187 30240 18199 30243
rect 19334 30240 19340 30252
rect 18187 30212 19340 30240
rect 18187 30209 18199 30212
rect 18141 30203 18199 30209
rect 19334 30200 19340 30212
rect 19392 30200 19398 30252
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 13173 30175 13231 30181
rect 13173 30172 13185 30175
rect 10735 30144 12020 30172
rect 12084 30144 12204 30172
rect 10735 30141 10747 30144
rect 10689 30135 10747 30141
rect 3108 30076 4752 30104
rect 9125 30107 9183 30113
rect 3108 30064 3114 30076
rect 9125 30073 9137 30107
rect 9171 30104 9183 30107
rect 9398 30104 9404 30116
rect 9171 30076 9404 30104
rect 9171 30073 9183 30076
rect 9125 30067 9183 30073
rect 9398 30064 9404 30076
rect 9456 30064 9462 30116
rect 2130 30036 2136 30048
rect 2091 30008 2136 30036
rect 2130 29996 2136 30008
rect 2188 29996 2194 30048
rect 2866 30036 2872 30048
rect 2827 30008 2872 30036
rect 2866 29996 2872 30008
rect 2924 29996 2930 30048
rect 7650 30036 7656 30048
rect 7611 30008 7656 30036
rect 7650 29996 7656 30008
rect 7708 29996 7714 30048
rect 8021 30039 8079 30045
rect 8021 30005 8033 30039
rect 8067 30036 8079 30039
rect 8938 30036 8944 30048
rect 8067 30008 8944 30036
rect 8067 30005 8079 30008
rect 8021 29999 8079 30005
rect 8938 29996 8944 30008
rect 8996 29996 9002 30048
rect 11701 30039 11759 30045
rect 11701 30005 11713 30039
rect 11747 30036 11759 30039
rect 11882 30036 11888 30048
rect 11747 30008 11888 30036
rect 11747 30005 11759 30008
rect 11701 29999 11759 30005
rect 11882 29996 11888 30008
rect 11940 29996 11946 30048
rect 11992 30036 12020 30144
rect 12176 30116 12204 30144
rect 12406 30144 13185 30172
rect 12158 30064 12164 30116
rect 12216 30104 12222 30116
rect 12406 30104 12434 30144
rect 13173 30141 13185 30144
rect 13219 30141 13231 30175
rect 17218 30172 17224 30184
rect 13173 30135 13231 30141
rect 13464 30144 17224 30172
rect 12216 30076 12434 30104
rect 12216 30064 12222 30076
rect 13464 30036 13492 30144
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 17957 30175 18015 30181
rect 17957 30172 17969 30175
rect 17512 30144 17969 30172
rect 17512 30116 17540 30144
rect 17957 30141 17969 30144
rect 18003 30172 18015 30175
rect 19150 30172 19156 30184
rect 18003 30144 19156 30172
rect 18003 30141 18015 30144
rect 17957 30135 18015 30141
rect 19150 30132 19156 30144
rect 19208 30172 19214 30184
rect 19628 30172 19656 30203
rect 20070 30200 20076 30252
rect 20128 30240 20134 30252
rect 20533 30243 20591 30249
rect 20533 30240 20545 30243
rect 20128 30212 20545 30240
rect 20128 30200 20134 30212
rect 20533 30209 20545 30212
rect 20579 30209 20591 30243
rect 22066 30240 22094 30280
rect 23106 30268 23112 30280
rect 23164 30268 23170 30320
rect 26050 30268 26056 30320
rect 26108 30308 26114 30320
rect 29748 30308 29776 30336
rect 30650 30317 30656 30320
rect 30627 30311 30656 30317
rect 26108 30280 29960 30308
rect 26108 30268 26114 30280
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 22066 30212 22385 30240
rect 20533 30203 20591 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 23014 30240 23020 30252
rect 22975 30212 23020 30240
rect 22373 30203 22431 30209
rect 23014 30200 23020 30212
rect 23072 30200 23078 30252
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23474 30240 23480 30252
rect 23247 30212 23480 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 23474 30200 23480 30212
rect 23532 30200 23538 30252
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30209 23903 30243
rect 23845 30203 23903 30209
rect 20257 30175 20315 30181
rect 20257 30172 20269 30175
rect 19208 30144 20269 30172
rect 19208 30132 19214 30144
rect 20257 30141 20269 30144
rect 20303 30141 20315 30175
rect 20257 30135 20315 30141
rect 22465 30175 22523 30181
rect 22465 30141 22477 30175
rect 22511 30172 22523 30175
rect 22738 30172 22744 30184
rect 22511 30144 22744 30172
rect 22511 30141 22523 30144
rect 22465 30135 22523 30141
rect 13541 30107 13599 30113
rect 13541 30073 13553 30107
rect 13587 30104 13599 30107
rect 13906 30104 13912 30116
rect 13587 30076 13912 30104
rect 13587 30073 13599 30076
rect 13541 30067 13599 30073
rect 13906 30064 13912 30076
rect 13964 30064 13970 30116
rect 14737 30107 14795 30113
rect 14737 30073 14749 30107
rect 14783 30104 14795 30107
rect 15838 30104 15844 30116
rect 14783 30076 15844 30104
rect 14783 30073 14795 30076
rect 14737 30067 14795 30073
rect 15838 30064 15844 30076
rect 15896 30104 15902 30116
rect 17494 30104 17500 30116
rect 15896 30076 17080 30104
rect 17455 30076 17500 30104
rect 15896 30064 15902 30076
rect 11992 30008 13492 30036
rect 13630 29996 13636 30048
rect 13688 30036 13694 30048
rect 14918 30036 14924 30048
rect 13688 30008 14924 30036
rect 13688 29996 13694 30008
rect 14918 29996 14924 30008
rect 14976 29996 14982 30048
rect 15102 29996 15108 30048
rect 15160 30036 15166 30048
rect 15381 30039 15439 30045
rect 15381 30036 15393 30039
rect 15160 30008 15393 30036
rect 15160 29996 15166 30008
rect 15381 30005 15393 30008
rect 15427 30005 15439 30039
rect 16942 30036 16948 30048
rect 16903 30008 16948 30036
rect 15381 29999 15439 30005
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 17052 30036 17080 30076
rect 17494 30064 17500 30076
rect 17552 30064 17558 30116
rect 17586 30064 17592 30116
rect 17644 30104 17650 30116
rect 19245 30107 19303 30113
rect 19245 30104 19257 30107
rect 17644 30076 19257 30104
rect 17644 30064 17650 30076
rect 19245 30073 19257 30076
rect 19291 30104 19303 30107
rect 19886 30104 19892 30116
rect 19291 30076 19892 30104
rect 19291 30073 19303 30076
rect 19245 30067 19303 30073
rect 19886 30064 19892 30076
rect 19944 30064 19950 30116
rect 19702 30036 19708 30048
rect 17052 30008 19708 30036
rect 19702 29996 19708 30008
rect 19760 29996 19766 30048
rect 19797 30039 19855 30045
rect 19797 30005 19809 30039
rect 19843 30036 19855 30039
rect 19978 30036 19984 30048
rect 19843 30008 19984 30036
rect 19843 30005 19855 30008
rect 19797 29999 19855 30005
rect 19978 29996 19984 30008
rect 20036 29996 20042 30048
rect 20272 30036 20300 30135
rect 22738 30132 22744 30144
rect 22796 30132 22802 30184
rect 22005 30107 22063 30113
rect 22005 30073 22017 30107
rect 22051 30104 22063 30107
rect 22370 30104 22376 30116
rect 22051 30076 22376 30104
rect 22051 30073 22063 30076
rect 22005 30067 22063 30073
rect 22370 30064 22376 30076
rect 22428 30064 22434 30116
rect 23860 30036 23888 30203
rect 24026 30200 24032 30252
rect 24084 30240 24090 30252
rect 25961 30243 26019 30249
rect 25961 30240 25973 30243
rect 24084 30212 25973 30240
rect 24084 30200 24090 30212
rect 25961 30209 25973 30212
rect 26007 30209 26019 30243
rect 25961 30203 26019 30209
rect 27709 30243 27767 30249
rect 27709 30209 27721 30243
rect 27755 30240 27767 30243
rect 27798 30240 27804 30252
rect 27755 30212 27804 30240
rect 27755 30209 27767 30212
rect 27709 30203 27767 30209
rect 27798 30200 27804 30212
rect 27856 30200 27862 30252
rect 27893 30243 27951 30249
rect 27893 30209 27905 30243
rect 27939 30240 27951 30243
rect 28626 30240 28632 30252
rect 27939 30212 28632 30240
rect 27939 30209 27951 30212
rect 27893 30203 27951 30209
rect 28626 30200 28632 30212
rect 28684 30200 28690 30252
rect 29661 30243 29719 30249
rect 29661 30209 29673 30243
rect 29707 30240 29719 30243
rect 29822 30240 29828 30252
rect 29707 30212 29828 30240
rect 29707 30209 29719 30212
rect 29661 30203 29719 30209
rect 29822 30200 29828 30212
rect 29880 30200 29886 30252
rect 29932 30249 29960 30280
rect 30627 30277 30639 30311
rect 30627 30271 30656 30277
rect 30650 30268 30656 30271
rect 30708 30268 30714 30320
rect 29917 30243 29975 30249
rect 29917 30209 29929 30243
rect 29963 30209 29975 30243
rect 29917 30203 29975 30209
rect 30006 30200 30012 30252
rect 30064 30240 30070 30252
rect 30502 30243 30560 30249
rect 30502 30240 30514 30243
rect 30064 30212 30514 30240
rect 30064 30200 30070 30212
rect 30502 30209 30514 30212
rect 30548 30209 30560 30243
rect 30502 30203 30560 30209
rect 31110 30200 31116 30252
rect 31168 30240 31174 30252
rect 31481 30243 31539 30249
rect 31481 30240 31493 30243
rect 31168 30212 31493 30240
rect 31168 30200 31174 30212
rect 31481 30209 31493 30212
rect 31527 30209 31539 30243
rect 31481 30203 31539 30209
rect 31570 30200 31576 30252
rect 31628 30240 31634 30252
rect 31757 30243 31815 30249
rect 31628 30212 31673 30240
rect 31628 30200 31634 30212
rect 31757 30209 31769 30243
rect 31803 30240 31815 30243
rect 32490 30240 32496 30252
rect 31803 30212 32496 30240
rect 31803 30209 31815 30212
rect 31757 30203 31815 30209
rect 32490 30200 32496 30212
rect 32548 30200 32554 30252
rect 32674 30240 32680 30252
rect 32635 30212 32680 30240
rect 32674 30200 32680 30212
rect 32732 30200 32738 30252
rect 37553 30243 37611 30249
rect 37553 30209 37565 30243
rect 37599 30240 37611 30243
rect 37642 30240 37648 30252
rect 37599 30212 37648 30240
rect 37599 30209 37611 30212
rect 37553 30203 37611 30209
rect 37642 30200 37648 30212
rect 37700 30200 37706 30252
rect 23937 30175 23995 30181
rect 23937 30141 23949 30175
rect 23983 30141 23995 30175
rect 23937 30135 23995 30141
rect 26053 30175 26111 30181
rect 26053 30141 26065 30175
rect 26099 30172 26111 30175
rect 26510 30172 26516 30184
rect 26099 30144 26516 30172
rect 26099 30141 26111 30144
rect 26053 30135 26111 30141
rect 20272 30008 23888 30036
rect 23952 30036 23980 30135
rect 26510 30132 26516 30144
rect 26568 30132 26574 30184
rect 28077 30175 28135 30181
rect 28077 30172 28089 30175
rect 27908 30144 28089 30172
rect 24213 30107 24271 30113
rect 24213 30073 24225 30107
rect 24259 30104 24271 30107
rect 24762 30104 24768 30116
rect 24259 30076 24768 30104
rect 24259 30073 24271 30076
rect 24213 30067 24271 30073
rect 24762 30064 24768 30076
rect 24820 30064 24826 30116
rect 26329 30107 26387 30113
rect 26329 30073 26341 30107
rect 26375 30104 26387 30107
rect 27522 30104 27528 30116
rect 26375 30076 27528 30104
rect 26375 30073 26387 30076
rect 26329 30067 26387 30073
rect 27522 30064 27528 30076
rect 27580 30064 27586 30116
rect 27614 30036 27620 30048
rect 23952 30008 27620 30036
rect 27614 29996 27620 30008
rect 27672 30036 27678 30048
rect 27908 30036 27936 30144
rect 28077 30141 28089 30144
rect 28123 30141 28135 30175
rect 28077 30135 28135 30141
rect 31021 30175 31079 30181
rect 31021 30141 31033 30175
rect 31067 30141 31079 30175
rect 31021 30135 31079 30141
rect 32585 30175 32643 30181
rect 32585 30141 32597 30175
rect 32631 30141 32643 30175
rect 32585 30135 32643 30141
rect 27672 30008 27936 30036
rect 28537 30039 28595 30045
rect 27672 29996 27678 30008
rect 28537 30005 28549 30039
rect 28583 30036 28595 30039
rect 28994 30036 29000 30048
rect 28583 30008 29000 30036
rect 28583 30005 28595 30008
rect 28537 29999 28595 30005
rect 28994 29996 29000 30008
rect 29052 29996 29058 30048
rect 29914 29996 29920 30048
rect 29972 30036 29978 30048
rect 30377 30039 30435 30045
rect 30377 30036 30389 30039
rect 29972 30008 30389 30036
rect 29972 29996 29978 30008
rect 30377 30005 30389 30008
rect 30423 30005 30435 30039
rect 30926 30036 30932 30048
rect 30887 30008 30932 30036
rect 30377 29999 30435 30005
rect 30926 29996 30932 30008
rect 30984 29996 30990 30048
rect 31036 30036 31064 30135
rect 31757 30107 31815 30113
rect 31757 30073 31769 30107
rect 31803 30104 31815 30107
rect 32600 30104 32628 30135
rect 31803 30076 32628 30104
rect 31803 30073 31815 30076
rect 31757 30067 31815 30073
rect 32401 30039 32459 30045
rect 32401 30036 32413 30039
rect 31036 30008 32413 30036
rect 32401 30005 32413 30008
rect 32447 30005 32459 30039
rect 32401 29999 32459 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 4433 29835 4491 29841
rect 4433 29801 4445 29835
rect 4479 29832 4491 29835
rect 4614 29832 4620 29844
rect 4479 29804 4620 29832
rect 4479 29801 4491 29804
rect 4433 29795 4491 29801
rect 4614 29792 4620 29804
rect 4672 29792 4678 29844
rect 5350 29832 5356 29844
rect 5311 29804 5356 29832
rect 5350 29792 5356 29804
rect 5408 29792 5414 29844
rect 10962 29792 10968 29844
rect 11020 29832 11026 29844
rect 11020 29804 11652 29832
rect 11020 29792 11026 29804
rect 9122 29764 9128 29776
rect 9083 29736 9128 29764
rect 9122 29724 9128 29736
rect 9180 29724 9186 29776
rect 11624 29764 11652 29804
rect 11974 29792 11980 29844
rect 12032 29832 12038 29844
rect 12069 29835 12127 29841
rect 12069 29832 12081 29835
rect 12032 29804 12081 29832
rect 12032 29792 12038 29804
rect 12069 29801 12081 29804
rect 12115 29801 12127 29835
rect 19794 29832 19800 29844
rect 12069 29795 12127 29801
rect 12176 29804 18092 29832
rect 19755 29804 19800 29832
rect 12176 29764 12204 29804
rect 14274 29764 14280 29776
rect 11624 29736 12204 29764
rect 14235 29736 14280 29764
rect 14274 29724 14280 29736
rect 14332 29724 14338 29776
rect 15286 29724 15292 29776
rect 15344 29764 15350 29776
rect 17494 29764 17500 29776
rect 15344 29736 17500 29764
rect 15344 29724 15350 29736
rect 17494 29724 17500 29736
rect 17552 29724 17558 29776
rect 17865 29767 17923 29773
rect 17865 29733 17877 29767
rect 17911 29764 17923 29767
rect 18064 29764 18092 29804
rect 19794 29792 19800 29804
rect 19852 29792 19858 29844
rect 20622 29832 20628 29844
rect 20583 29804 20628 29832
rect 20622 29792 20628 29804
rect 20680 29792 20686 29844
rect 21821 29835 21879 29841
rect 21821 29801 21833 29835
rect 21867 29832 21879 29835
rect 22094 29832 22100 29844
rect 21867 29804 22100 29832
rect 21867 29801 21879 29804
rect 21821 29795 21879 29801
rect 22094 29792 22100 29804
rect 22152 29792 22158 29844
rect 24854 29792 24860 29844
rect 24912 29832 24918 29844
rect 25041 29835 25099 29841
rect 25041 29832 25053 29835
rect 24912 29804 25053 29832
rect 24912 29792 24918 29804
rect 25041 29801 25053 29804
rect 25087 29801 25099 29835
rect 25041 29795 25099 29801
rect 26234 29792 26240 29844
rect 26292 29832 26298 29844
rect 28445 29835 28503 29841
rect 28445 29832 28457 29835
rect 26292 29804 28457 29832
rect 26292 29792 26298 29804
rect 28445 29801 28457 29804
rect 28491 29801 28503 29835
rect 28626 29832 28632 29844
rect 28587 29804 28632 29832
rect 28445 29795 28503 29801
rect 28626 29792 28632 29804
rect 28684 29792 28690 29844
rect 29822 29792 29828 29844
rect 29880 29832 29886 29844
rect 29917 29835 29975 29841
rect 29917 29832 29929 29835
rect 29880 29804 29929 29832
rect 29880 29792 29886 29804
rect 29917 29801 29929 29804
rect 29963 29801 29975 29835
rect 30558 29832 30564 29844
rect 30519 29804 30564 29832
rect 29917 29795 29975 29801
rect 30558 29792 30564 29804
rect 30616 29792 30622 29844
rect 33594 29832 33600 29844
rect 31726 29804 33600 29832
rect 31726 29764 31754 29804
rect 33594 29792 33600 29804
rect 33652 29832 33658 29844
rect 38378 29832 38384 29844
rect 33652 29804 38384 29832
rect 33652 29792 33658 29804
rect 38378 29792 38384 29804
rect 38436 29792 38442 29844
rect 17911 29736 18000 29764
rect 18064 29736 31754 29764
rect 17911 29733 17923 29736
rect 17865 29727 17923 29733
rect 2958 29656 2964 29708
rect 3016 29696 3022 29708
rect 3421 29699 3479 29705
rect 3421 29696 3433 29699
rect 3016 29668 3433 29696
rect 3016 29656 3022 29668
rect 3421 29665 3433 29668
rect 3467 29665 3479 29699
rect 10134 29696 10140 29708
rect 3421 29659 3479 29665
rect 5092 29668 10140 29696
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29628 4583 29631
rect 4614 29628 4620 29640
rect 4571 29600 4620 29628
rect 4571 29597 4583 29600
rect 4525 29591 4583 29597
rect 4614 29588 4620 29600
rect 4672 29588 4678 29640
rect 1578 29560 1584 29572
rect 1539 29532 1584 29560
rect 1578 29520 1584 29532
rect 1636 29520 1642 29572
rect 3234 29560 3240 29572
rect 3195 29532 3240 29560
rect 3234 29520 3240 29532
rect 3292 29520 3298 29572
rect 5092 29569 5120 29668
rect 10134 29656 10140 29668
rect 10192 29656 10198 29708
rect 15654 29656 15660 29708
rect 15712 29696 15718 29708
rect 17972 29696 18000 29736
rect 18598 29696 18604 29708
rect 15712 29668 17908 29696
rect 17972 29668 18604 29696
rect 15712 29656 15718 29668
rect 7650 29588 7656 29640
rect 7708 29628 7714 29640
rect 9309 29631 9367 29637
rect 9309 29628 9321 29631
rect 7708 29600 9321 29628
rect 7708 29588 7714 29600
rect 9309 29597 9321 29600
rect 9355 29597 9367 29631
rect 9309 29591 9367 29597
rect 9401 29631 9459 29637
rect 9401 29597 9413 29631
rect 9447 29628 9459 29631
rect 9582 29628 9588 29640
rect 9447 29600 9588 29628
rect 9447 29597 9459 29600
rect 9401 29591 9459 29597
rect 9582 29588 9588 29600
rect 9640 29588 9646 29640
rect 10042 29628 10048 29640
rect 10003 29600 10048 29628
rect 10042 29588 10048 29600
rect 10100 29588 10106 29640
rect 10689 29631 10747 29637
rect 10689 29597 10701 29631
rect 10735 29628 10747 29631
rect 12434 29628 12440 29640
rect 10735 29600 12440 29628
rect 10735 29597 10747 29600
rect 10689 29591 10747 29597
rect 12434 29588 12440 29600
rect 12492 29588 12498 29640
rect 12529 29631 12587 29637
rect 12529 29597 12541 29631
rect 12575 29597 12587 29631
rect 12529 29591 12587 29597
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29628 13507 29631
rect 13630 29628 13636 29640
rect 13495 29600 13636 29628
rect 13495 29597 13507 29600
rect 13449 29591 13507 29597
rect 5077 29563 5135 29569
rect 5077 29529 5089 29563
rect 5123 29529 5135 29563
rect 5077 29523 5135 29529
rect 2958 29452 2964 29504
rect 3016 29492 3022 29504
rect 5092 29492 5120 29523
rect 9030 29520 9036 29572
rect 9088 29560 9094 29572
rect 9125 29563 9183 29569
rect 9125 29560 9137 29563
rect 9088 29532 9137 29560
rect 9088 29520 9094 29532
rect 9125 29529 9137 29532
rect 9171 29529 9183 29563
rect 10934 29563 10992 29569
rect 10934 29560 10946 29563
rect 9125 29523 9183 29529
rect 10244 29532 10946 29560
rect 10244 29501 10272 29532
rect 10934 29529 10946 29532
rect 10980 29529 10992 29563
rect 10934 29523 10992 29529
rect 11974 29520 11980 29572
rect 12032 29560 12038 29572
rect 12544 29560 12572 29591
rect 13630 29588 13636 29600
rect 13688 29588 13694 29640
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 14274 29628 14280 29640
rect 13771 29600 14280 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 14458 29637 14464 29640
rect 14436 29631 14464 29637
rect 14436 29597 14448 29631
rect 14436 29591 14464 29597
rect 14458 29588 14464 29591
rect 14516 29588 14522 29640
rect 14734 29588 14740 29640
rect 14792 29637 14798 29640
rect 14792 29631 14831 29637
rect 14819 29597 14831 29631
rect 14792 29591 14831 29597
rect 14792 29588 14798 29591
rect 14918 29588 14924 29640
rect 14976 29628 14982 29640
rect 14976 29600 15021 29628
rect 14976 29588 14982 29600
rect 15378 29588 15384 29640
rect 15436 29628 15442 29640
rect 15565 29631 15623 29637
rect 15565 29628 15577 29631
rect 15436 29600 15577 29628
rect 15436 29588 15442 29600
rect 15565 29597 15577 29600
rect 15611 29597 15623 29631
rect 15565 29591 15623 29597
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29628 15807 29631
rect 17126 29628 17132 29640
rect 15795 29600 17132 29628
rect 15795 29597 15807 29600
rect 15749 29591 15807 29597
rect 17126 29588 17132 29600
rect 17184 29588 17190 29640
rect 17405 29631 17463 29637
rect 17405 29597 17417 29631
rect 17451 29628 17463 29631
rect 17770 29628 17776 29640
rect 17451 29600 17776 29628
rect 17451 29597 17463 29600
rect 17405 29591 17463 29597
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 17880 29628 17908 29668
rect 18598 29656 18604 29668
rect 18656 29656 18662 29708
rect 19613 29699 19671 29705
rect 19613 29665 19625 29699
rect 19659 29696 19671 29699
rect 23014 29696 23020 29708
rect 19659 29668 23020 29696
rect 19659 29665 19671 29668
rect 19613 29659 19671 29665
rect 19628 29628 19656 29659
rect 23014 29656 23020 29668
rect 23072 29656 23078 29708
rect 24670 29696 24676 29708
rect 24631 29668 24676 29696
rect 24670 29656 24676 29668
rect 24728 29656 24734 29708
rect 26694 29696 26700 29708
rect 26655 29668 26700 29696
rect 26694 29656 26700 29668
rect 26752 29656 26758 29708
rect 30926 29656 30932 29708
rect 30984 29696 30990 29708
rect 31113 29699 31171 29705
rect 31113 29696 31125 29699
rect 30984 29668 31125 29696
rect 30984 29656 30990 29668
rect 31113 29665 31125 29668
rect 31159 29665 31171 29699
rect 37182 29696 37188 29708
rect 37143 29668 37188 29696
rect 31113 29659 31171 29665
rect 37182 29656 37188 29668
rect 37240 29656 37246 29708
rect 17880 29600 19656 29628
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 13354 29560 13360 29572
rect 12032 29532 12572 29560
rect 12728 29532 13360 29560
rect 12032 29520 12038 29532
rect 12728 29504 12756 29532
rect 13354 29520 13360 29532
rect 13412 29560 13418 29572
rect 14553 29563 14611 29569
rect 14553 29560 14565 29563
rect 13412 29532 14565 29560
rect 13412 29520 13418 29532
rect 14553 29529 14565 29532
rect 14599 29529 14611 29563
rect 14553 29523 14611 29529
rect 14645 29563 14703 29569
rect 14645 29529 14657 29563
rect 14691 29529 14703 29563
rect 14645 29523 14703 29529
rect 3016 29464 5120 29492
rect 10229 29495 10287 29501
rect 3016 29452 3022 29464
rect 10229 29461 10241 29495
rect 10275 29461 10287 29495
rect 10229 29455 10287 29461
rect 12621 29495 12679 29501
rect 12621 29461 12633 29495
rect 12667 29492 12679 29495
rect 12710 29492 12716 29504
rect 12667 29464 12716 29492
rect 12667 29461 12679 29464
rect 12621 29455 12679 29461
rect 12710 29452 12716 29464
rect 12768 29452 12774 29504
rect 13262 29492 13268 29504
rect 13223 29464 13268 29492
rect 13262 29452 13268 29464
rect 13320 29452 13326 29504
rect 13633 29495 13691 29501
rect 13633 29461 13645 29495
rect 13679 29492 13691 29495
rect 13814 29492 13820 29504
rect 13679 29464 13820 29492
rect 13679 29461 13691 29464
rect 13633 29455 13691 29461
rect 13814 29452 13820 29464
rect 13872 29492 13878 29504
rect 14660 29492 14688 29523
rect 16850 29520 16856 29572
rect 16908 29560 16914 29572
rect 17313 29563 17371 29569
rect 17313 29560 17325 29563
rect 16908 29532 17325 29560
rect 16908 29520 16914 29532
rect 17313 29529 17325 29532
rect 17359 29529 17371 29563
rect 17313 29523 17371 29529
rect 17865 29563 17923 29569
rect 17865 29529 17877 29563
rect 17911 29560 17923 29563
rect 18782 29560 18788 29572
rect 17911 29532 18788 29560
rect 17911 29529 17923 29532
rect 17865 29523 17923 29529
rect 18782 29520 18788 29532
rect 18840 29520 18846 29572
rect 19518 29520 19524 29572
rect 19576 29560 19582 29572
rect 19720 29560 19748 29591
rect 19886 29588 19892 29640
rect 19944 29588 19950 29640
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29628 20039 29631
rect 20070 29628 20076 29640
rect 20027 29600 20076 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 20438 29588 20444 29640
rect 20496 29628 20502 29640
rect 20625 29631 20683 29637
rect 20625 29628 20637 29631
rect 20496 29600 20637 29628
rect 20496 29588 20502 29600
rect 20625 29597 20637 29600
rect 20671 29597 20683 29631
rect 20806 29628 20812 29640
rect 20767 29600 20812 29628
rect 20625 29591 20683 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 20898 29588 20904 29640
rect 20956 29628 20962 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 20956 29600 24777 29628
rect 20956 29588 20962 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 26510 29628 26516 29640
rect 26471 29600 26516 29628
rect 24765 29591 24823 29597
rect 26510 29588 26516 29600
rect 26568 29588 26574 29640
rect 29730 29628 29736 29640
rect 29691 29600 29736 29628
rect 29730 29588 29736 29600
rect 29788 29588 29794 29640
rect 29914 29628 29920 29640
rect 29875 29600 29920 29628
rect 29914 29588 29920 29600
rect 29972 29588 29978 29640
rect 30742 29631 30800 29637
rect 30742 29597 30754 29631
rect 30788 29628 30800 29631
rect 31018 29628 31024 29640
rect 30788 29600 31024 29628
rect 30788 29597 30800 29600
rect 30742 29591 30800 29597
rect 31018 29588 31024 29600
rect 31076 29588 31082 29640
rect 31205 29631 31263 29637
rect 31205 29597 31217 29631
rect 31251 29628 31263 29631
rect 32125 29631 32183 29637
rect 32125 29628 32137 29631
rect 31251 29600 32137 29628
rect 31251 29597 31263 29600
rect 31205 29591 31263 29597
rect 32125 29597 32137 29600
rect 32171 29597 32183 29631
rect 32125 29591 32183 29597
rect 38286 29588 38292 29640
rect 38344 29628 38350 29640
rect 38344 29600 38389 29628
rect 38344 29588 38350 29600
rect 19576 29532 19748 29560
rect 19904 29560 19932 29588
rect 22005 29563 22063 29569
rect 22005 29560 22017 29563
rect 19904 29532 22017 29560
rect 19576 29520 19582 29532
rect 22005 29529 22017 29532
rect 22051 29529 22063 29563
rect 22005 29523 22063 29529
rect 22189 29563 22247 29569
rect 22189 29529 22201 29563
rect 22235 29560 22247 29563
rect 23474 29560 23480 29572
rect 22235 29532 23480 29560
rect 22235 29529 22247 29532
rect 22189 29523 22247 29529
rect 23474 29520 23480 29532
rect 23532 29560 23538 29572
rect 23750 29560 23756 29572
rect 23532 29532 23756 29560
rect 23532 29520 23538 29532
rect 23750 29520 23756 29532
rect 23808 29520 23814 29572
rect 27246 29560 27252 29572
rect 27159 29532 27252 29560
rect 27246 29520 27252 29532
rect 27304 29560 27310 29572
rect 27890 29560 27896 29572
rect 27304 29532 27896 29560
rect 27304 29520 27310 29532
rect 27890 29520 27896 29532
rect 27948 29520 27954 29572
rect 28813 29563 28871 29569
rect 28813 29529 28825 29563
rect 28859 29560 28871 29563
rect 28994 29560 29000 29572
rect 28859 29532 29000 29560
rect 28859 29529 28871 29532
rect 28813 29523 28871 29529
rect 28994 29520 29000 29532
rect 29052 29520 29058 29572
rect 32306 29560 32312 29572
rect 32267 29532 32312 29560
rect 32306 29520 32312 29532
rect 32364 29520 32370 29572
rect 32490 29560 32496 29572
rect 32451 29532 32496 29560
rect 32490 29520 32496 29532
rect 32548 29520 32554 29572
rect 38102 29560 38108 29572
rect 38063 29532 38108 29560
rect 38102 29520 38108 29532
rect 38160 29520 38166 29572
rect 13872 29464 14688 29492
rect 15381 29495 15439 29501
rect 13872 29452 13878 29464
rect 15381 29461 15393 29495
rect 15427 29492 15439 29495
rect 15562 29492 15568 29504
rect 15427 29464 15568 29492
rect 15427 29461 15439 29464
rect 15381 29455 15439 29461
rect 15562 29452 15568 29464
rect 15620 29452 15626 29504
rect 17129 29495 17187 29501
rect 17129 29461 17141 29495
rect 17175 29492 17187 29495
rect 19426 29492 19432 29504
rect 17175 29464 19432 29492
rect 17175 29461 17187 29464
rect 17129 29455 17187 29461
rect 19426 29452 19432 29464
rect 19484 29452 19490 29504
rect 19889 29495 19947 29501
rect 19889 29461 19901 29495
rect 19935 29492 19947 29495
rect 20070 29492 20076 29504
rect 19935 29464 20076 29492
rect 19935 29461 19947 29464
rect 19889 29455 19947 29461
rect 20070 29452 20076 29464
rect 20128 29452 20134 29504
rect 27338 29492 27344 29504
rect 27299 29464 27344 29492
rect 27338 29452 27344 29464
rect 27396 29452 27402 29504
rect 28613 29495 28671 29501
rect 28613 29461 28625 29495
rect 28659 29492 28671 29495
rect 29086 29492 29092 29504
rect 28659 29464 29092 29492
rect 28659 29461 28671 29464
rect 28613 29455 28671 29461
rect 29086 29452 29092 29464
rect 29144 29452 29150 29504
rect 30650 29452 30656 29504
rect 30708 29492 30714 29504
rect 30745 29495 30803 29501
rect 30745 29492 30757 29495
rect 30708 29464 30757 29492
rect 30708 29452 30714 29464
rect 30745 29461 30757 29464
rect 30791 29461 30803 29495
rect 30745 29455 30803 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 10042 29248 10048 29300
rect 10100 29288 10106 29300
rect 11701 29291 11759 29297
rect 11701 29288 11713 29291
rect 10100 29260 11713 29288
rect 10100 29248 10106 29260
rect 11701 29257 11713 29260
rect 11747 29257 11759 29291
rect 11882 29288 11888 29300
rect 11843 29260 11888 29288
rect 11701 29251 11759 29257
rect 11882 29248 11888 29260
rect 11940 29248 11946 29300
rect 12434 29248 12440 29300
rect 12492 29288 12498 29300
rect 16758 29288 16764 29300
rect 12492 29260 16764 29288
rect 12492 29248 12498 29260
rect 16758 29248 16764 29260
rect 16816 29288 16822 29300
rect 16942 29288 16948 29300
rect 16816 29260 16948 29288
rect 16816 29248 16822 29260
rect 16942 29248 16948 29260
rect 17000 29248 17006 29300
rect 17218 29248 17224 29300
rect 17276 29288 17282 29300
rect 31573 29291 31631 29297
rect 17276 29260 31524 29288
rect 17276 29248 17282 29260
rect 18316 29223 18374 29229
rect 6886 29192 17264 29220
rect 2130 29152 2136 29164
rect 2091 29124 2136 29152
rect 2130 29112 2136 29124
rect 2188 29112 2194 29164
rect 4801 29155 4859 29161
rect 4801 29121 4813 29155
rect 4847 29152 4859 29155
rect 5350 29152 5356 29164
rect 4847 29124 5356 29152
rect 4847 29121 4859 29124
rect 4801 29115 4859 29121
rect 5350 29112 5356 29124
rect 5408 29112 5414 29164
rect 2317 29087 2375 29093
rect 2317 29053 2329 29087
rect 2363 29084 2375 29087
rect 2774 29084 2780 29096
rect 2363 29056 2780 29084
rect 2363 29053 2375 29056
rect 2317 29047 2375 29053
rect 2774 29044 2780 29056
rect 2832 29044 2838 29096
rect 2866 29044 2872 29096
rect 2924 29084 2930 29096
rect 2924 29056 2969 29084
rect 2924 29044 2930 29056
rect 4614 28976 4620 29028
rect 4672 29016 4678 29028
rect 6886 29016 6914 29192
rect 8205 29155 8263 29161
rect 8205 29121 8217 29155
rect 8251 29152 8263 29155
rect 8662 29152 8668 29164
rect 8251 29124 8668 29152
rect 8251 29121 8263 29124
rect 8205 29115 8263 29121
rect 8662 29112 8668 29124
rect 8720 29112 8726 29164
rect 10134 29112 10140 29164
rect 10192 29152 10198 29164
rect 10413 29155 10471 29161
rect 10413 29152 10425 29155
rect 10192 29124 10425 29152
rect 10192 29112 10198 29124
rect 10413 29121 10425 29124
rect 10459 29121 10471 29155
rect 10962 29152 10968 29164
rect 10923 29124 10968 29152
rect 10413 29115 10471 29121
rect 10962 29112 10968 29124
rect 11020 29112 11026 29164
rect 11790 29112 11796 29164
rect 11848 29152 11854 29164
rect 12253 29155 12311 29161
rect 12253 29152 12265 29155
rect 11848 29124 12265 29152
rect 11848 29112 11854 29124
rect 12253 29121 12265 29124
rect 12299 29121 12311 29155
rect 13357 29155 13415 29161
rect 13357 29152 13369 29155
rect 12253 29115 12311 29121
rect 12406 29124 13369 29152
rect 8113 29087 8171 29093
rect 8113 29053 8125 29087
rect 8159 29053 8171 29087
rect 8113 29047 8171 29053
rect 4672 28988 6914 29016
rect 8128 29016 8156 29047
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10980 29084 11008 29112
rect 9732 29056 11008 29084
rect 9732 29044 9738 29056
rect 12158 29044 12164 29096
rect 12216 29084 12222 29096
rect 12406 29084 12434 29124
rect 13357 29121 13369 29124
rect 13403 29121 13415 29155
rect 13357 29115 13415 29121
rect 15013 29155 15071 29161
rect 15013 29121 15025 29155
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 13814 29084 13820 29096
rect 12216 29056 12434 29084
rect 13775 29056 13820 29084
rect 12216 29044 12222 29056
rect 13814 29044 13820 29056
rect 13872 29044 13878 29096
rect 14274 29044 14280 29096
rect 14332 29084 14338 29096
rect 14553 29087 14611 29093
rect 14553 29084 14565 29087
rect 14332 29056 14565 29084
rect 14332 29044 14338 29056
rect 14553 29053 14565 29056
rect 14599 29084 14611 29087
rect 14734 29084 14740 29096
rect 14599 29056 14740 29084
rect 14599 29053 14611 29056
rect 14553 29047 14611 29053
rect 14734 29044 14740 29056
rect 14792 29044 14798 29096
rect 15028 29084 15056 29115
rect 15102 29112 15108 29164
rect 15160 29152 15166 29164
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 15160 29124 16865 29152
rect 15160 29112 15166 29124
rect 16853 29121 16865 29124
rect 16899 29121 16911 29155
rect 16853 29115 16911 29121
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29152 17095 29155
rect 17126 29152 17132 29164
rect 17083 29124 17132 29152
rect 17083 29121 17095 29124
rect 17037 29115 17095 29121
rect 17126 29112 17132 29124
rect 17184 29112 17190 29164
rect 17236 29152 17264 29192
rect 18316 29189 18328 29223
rect 18362 29220 18374 29223
rect 18690 29220 18696 29232
rect 18362 29192 18696 29220
rect 18362 29189 18374 29192
rect 18316 29183 18374 29189
rect 18690 29180 18696 29192
rect 18748 29180 18754 29232
rect 18782 29180 18788 29232
rect 18840 29220 18846 29232
rect 24026 29220 24032 29232
rect 18840 29192 24032 29220
rect 18840 29180 18846 29192
rect 24026 29180 24032 29192
rect 24084 29180 24090 29232
rect 25133 29223 25191 29229
rect 25133 29189 25145 29223
rect 25179 29220 25191 29223
rect 25958 29220 25964 29232
rect 25179 29192 25964 29220
rect 25179 29189 25191 29192
rect 25133 29183 25191 29189
rect 25958 29180 25964 29192
rect 26016 29180 26022 29232
rect 30745 29223 30803 29229
rect 30745 29189 30757 29223
rect 30791 29220 30803 29223
rect 31389 29223 31447 29229
rect 31389 29220 31401 29223
rect 30791 29192 31401 29220
rect 30791 29189 30803 29192
rect 30745 29183 30803 29189
rect 31389 29189 31401 29192
rect 31435 29189 31447 29223
rect 31496 29220 31524 29260
rect 31573 29257 31585 29291
rect 31619 29288 31631 29291
rect 32674 29288 32680 29300
rect 31619 29260 32680 29288
rect 31619 29257 31631 29260
rect 31573 29251 31631 29257
rect 32674 29248 32680 29260
rect 32732 29248 32738 29300
rect 37642 29220 37648 29232
rect 31496 29192 37648 29220
rect 31389 29183 31447 29189
rect 37642 29180 37648 29192
rect 37700 29180 37706 29232
rect 20993 29155 21051 29161
rect 17236 29124 19104 29152
rect 15654 29084 15660 29096
rect 15028 29056 15660 29084
rect 15654 29044 15660 29056
rect 15712 29084 15718 29096
rect 15933 29087 15991 29093
rect 15933 29084 15945 29087
rect 15712 29056 15945 29084
rect 15712 29044 15718 29056
rect 15933 29053 15945 29056
rect 15979 29053 15991 29087
rect 15933 29047 15991 29053
rect 16942 29044 16948 29096
rect 17000 29084 17006 29096
rect 18049 29087 18107 29093
rect 18049 29084 18061 29087
rect 17000 29056 18061 29084
rect 17000 29044 17006 29056
rect 18049 29053 18061 29056
rect 18095 29053 18107 29087
rect 19076 29084 19104 29124
rect 20993 29121 21005 29155
rect 21039 29152 21051 29155
rect 21082 29152 21088 29164
rect 21039 29124 21088 29152
rect 21039 29121 21051 29124
rect 20993 29115 21051 29121
rect 21082 29112 21088 29124
rect 21140 29112 21146 29164
rect 21174 29112 21180 29164
rect 21232 29152 21238 29164
rect 23382 29152 23388 29164
rect 21232 29124 21277 29152
rect 23343 29124 23388 29152
rect 21232 29112 21238 29124
rect 23382 29112 23388 29124
rect 23440 29112 23446 29164
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29121 26479 29155
rect 26421 29115 26479 29121
rect 25406 29084 25412 29096
rect 19076 29056 25412 29084
rect 18049 29047 18107 29053
rect 15286 29016 15292 29028
rect 8128 28988 15292 29016
rect 4672 28976 4678 28988
rect 15286 28976 15292 28988
rect 15344 28976 15350 29028
rect 15470 29016 15476 29028
rect 15431 28988 15476 29016
rect 15470 28976 15476 28988
rect 15528 28976 15534 29028
rect 15562 28976 15568 29028
rect 15620 29016 15626 29028
rect 15620 28988 15665 29016
rect 15620 28976 15626 28988
rect 15746 28976 15752 29028
rect 15804 29016 15810 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 15804 28988 16865 29016
rect 15804 28976 15810 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16853 28979 16911 28985
rect 4706 28948 4712 28960
rect 4667 28920 4712 28948
rect 4706 28908 4712 28920
rect 4764 28908 4770 28960
rect 7834 28948 7840 28960
rect 7795 28920 7840 28948
rect 7834 28908 7840 28920
rect 7892 28908 7898 28960
rect 11882 28948 11888 28960
rect 11843 28920 11888 28948
rect 11882 28908 11888 28920
rect 11940 28908 11946 28960
rect 13633 28951 13691 28957
rect 13633 28917 13645 28951
rect 13679 28948 13691 28951
rect 13906 28948 13912 28960
rect 13679 28920 13912 28948
rect 13679 28917 13691 28920
rect 13633 28911 13691 28917
rect 13906 28908 13912 28920
rect 13964 28908 13970 28960
rect 14921 28951 14979 28957
rect 14921 28917 14933 28951
rect 14967 28948 14979 28951
rect 15378 28948 15384 28960
rect 14967 28920 15384 28948
rect 14967 28917 14979 28920
rect 14921 28911 14979 28917
rect 15378 28908 15384 28920
rect 15436 28908 15442 28960
rect 18064 28948 18092 29047
rect 25406 29044 25412 29056
rect 25464 29044 25470 29096
rect 19150 28976 19156 29028
rect 19208 29016 19214 29028
rect 19429 29019 19487 29025
rect 19429 29016 19441 29019
rect 19208 28988 19441 29016
rect 19208 28976 19214 28988
rect 19429 28985 19441 28988
rect 19475 28985 19487 29019
rect 19429 28979 19487 28985
rect 26237 29019 26295 29025
rect 26237 28985 26249 29019
rect 26283 29016 26295 29019
rect 26326 29016 26332 29028
rect 26283 28988 26332 29016
rect 26283 28985 26295 28988
rect 26237 28979 26295 28985
rect 26326 28976 26332 28988
rect 26384 28976 26390 29028
rect 26436 28960 26464 29115
rect 30006 29112 30012 29164
rect 30064 29152 30070 29164
rect 30561 29155 30619 29161
rect 30561 29152 30573 29155
rect 30064 29124 30573 29152
rect 30064 29112 30070 29124
rect 30561 29121 30573 29124
rect 30607 29121 30619 29155
rect 30561 29115 30619 29121
rect 31018 29112 31024 29164
rect 31076 29152 31082 29164
rect 31205 29155 31263 29161
rect 31205 29152 31217 29155
rect 31076 29124 31217 29152
rect 31076 29112 31082 29124
rect 31205 29121 31217 29124
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 37829 29155 37887 29161
rect 37829 29121 37841 29155
rect 37875 29152 37887 29155
rect 38286 29152 38292 29164
rect 37875 29124 38292 29152
rect 37875 29121 37887 29124
rect 37829 29115 37887 29121
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 30374 29084 30380 29096
rect 30287 29056 30380 29084
rect 30374 29044 30380 29056
rect 30432 29084 30438 29096
rect 31570 29084 31576 29096
rect 30432 29056 31576 29084
rect 30432 29044 30438 29056
rect 31570 29044 31576 29056
rect 31628 29044 31634 29096
rect 18414 28948 18420 28960
rect 18064 28920 18420 28948
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 21085 28951 21143 28957
rect 21085 28917 21097 28951
rect 21131 28948 21143 28951
rect 21174 28948 21180 28960
rect 21131 28920 21180 28948
rect 21131 28917 21143 28920
rect 21085 28911 21143 28917
rect 21174 28908 21180 28920
rect 21232 28908 21238 28960
rect 26418 28908 26424 28960
rect 26476 28948 26482 28960
rect 31386 28948 31392 28960
rect 26476 28920 31392 28948
rect 26476 28908 26482 28920
rect 31386 28908 31392 28920
rect 31444 28908 31450 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 2774 28744 2780 28756
rect 2735 28716 2780 28744
rect 2774 28704 2780 28716
rect 2832 28704 2838 28756
rect 11790 28744 11796 28756
rect 11751 28716 11796 28744
rect 11790 28704 11796 28716
rect 11848 28704 11854 28756
rect 11977 28747 12035 28753
rect 11977 28713 11989 28747
rect 12023 28744 12035 28747
rect 12158 28744 12164 28756
rect 12023 28716 12164 28744
rect 12023 28713 12035 28716
rect 11977 28707 12035 28713
rect 12158 28704 12164 28716
rect 12216 28704 12222 28756
rect 16942 28744 16948 28756
rect 16903 28716 16948 28744
rect 16942 28704 16948 28716
rect 17000 28704 17006 28756
rect 26510 28704 26516 28756
rect 26568 28744 26574 28756
rect 26605 28747 26663 28753
rect 26605 28744 26617 28747
rect 26568 28716 26617 28744
rect 26568 28704 26574 28716
rect 26605 28713 26617 28716
rect 26651 28713 26663 28747
rect 28166 28744 28172 28756
rect 28127 28716 28172 28744
rect 26605 28707 26663 28713
rect 28166 28704 28172 28716
rect 28224 28704 28230 28756
rect 38102 28704 38108 28756
rect 38160 28744 38166 28756
rect 38197 28747 38255 28753
rect 38197 28744 38209 28747
rect 38160 28716 38209 28744
rect 38160 28704 38166 28716
rect 38197 28713 38209 28716
rect 38243 28713 38255 28747
rect 38197 28707 38255 28713
rect 20073 28679 20131 28685
rect 20073 28645 20085 28679
rect 20119 28676 20131 28679
rect 20254 28676 20260 28688
rect 20119 28648 20260 28676
rect 20119 28645 20131 28648
rect 20073 28639 20131 28645
rect 20254 28636 20260 28648
rect 20312 28636 20318 28688
rect 31205 28679 31263 28685
rect 31205 28645 31217 28679
rect 31251 28676 31263 28679
rect 31570 28676 31576 28688
rect 31251 28648 31576 28676
rect 31251 28645 31263 28648
rect 31205 28639 31263 28645
rect 31570 28636 31576 28648
rect 31628 28636 31634 28688
rect 4433 28611 4491 28617
rect 4433 28577 4445 28611
rect 4479 28608 4491 28611
rect 4706 28608 4712 28620
rect 4479 28580 4712 28608
rect 4479 28577 4491 28580
rect 4433 28571 4491 28577
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 5626 28608 5632 28620
rect 5587 28580 5632 28608
rect 5626 28568 5632 28580
rect 5684 28568 5690 28620
rect 7834 28568 7840 28620
rect 7892 28608 7898 28620
rect 8113 28611 8171 28617
rect 8113 28608 8125 28611
rect 7892 28580 8125 28608
rect 7892 28568 7898 28580
rect 8113 28577 8125 28580
rect 8159 28577 8171 28611
rect 8113 28571 8171 28577
rect 11882 28568 11888 28620
rect 11940 28608 11946 28620
rect 17310 28608 17316 28620
rect 11940 28580 17316 28608
rect 11940 28568 11946 28580
rect 17310 28568 17316 28580
rect 17368 28608 17374 28620
rect 21266 28608 21272 28620
rect 17368 28580 18552 28608
rect 17368 28568 17374 28580
rect 1854 28500 1860 28552
rect 1912 28540 1918 28552
rect 1949 28543 2007 28549
rect 1949 28540 1961 28543
rect 1912 28512 1961 28540
rect 1912 28500 1918 28512
rect 1949 28509 1961 28512
rect 1995 28509 2007 28543
rect 1949 28503 2007 28509
rect 2869 28543 2927 28549
rect 2869 28509 2881 28543
rect 2915 28540 2927 28543
rect 2958 28540 2964 28552
rect 2915 28512 2964 28540
rect 2915 28509 2927 28512
rect 2869 28503 2927 28509
rect 2958 28500 2964 28512
rect 3016 28500 3022 28552
rect 4246 28540 4252 28552
rect 4207 28512 4252 28540
rect 4246 28500 4252 28512
rect 4304 28500 4310 28552
rect 8205 28543 8263 28549
rect 8205 28509 8217 28543
rect 8251 28540 8263 28543
rect 9122 28540 9128 28552
rect 8251 28512 9128 28540
rect 8251 28509 8263 28512
rect 8205 28503 8263 28509
rect 9122 28500 9128 28512
rect 9180 28500 9186 28552
rect 11974 28500 11980 28552
rect 12032 28500 12038 28552
rect 15657 28543 15715 28549
rect 15657 28509 15669 28543
rect 15703 28540 15715 28543
rect 17402 28540 17408 28552
rect 15703 28512 17408 28540
rect 15703 28509 15715 28512
rect 15657 28503 15715 28509
rect 17402 28500 17408 28512
rect 17460 28500 17466 28552
rect 18524 28549 18552 28580
rect 20364 28580 21272 28608
rect 20364 28549 20392 28580
rect 21266 28568 21272 28580
rect 21324 28568 21330 28620
rect 27614 28568 27620 28620
rect 27672 28608 27678 28620
rect 28261 28611 28319 28617
rect 28261 28608 28273 28611
rect 27672 28580 28273 28608
rect 27672 28568 27678 28580
rect 28261 28577 28273 28580
rect 28307 28608 28319 28611
rect 30006 28608 30012 28620
rect 28307 28580 30012 28608
rect 28307 28577 28319 28580
rect 28261 28571 28319 28577
rect 30006 28568 30012 28580
rect 30064 28568 30070 28620
rect 37645 28611 37703 28617
rect 37645 28577 37657 28611
rect 37691 28608 37703 28611
rect 37734 28608 37740 28620
rect 37691 28580 37740 28608
rect 37691 28577 37703 28580
rect 37645 28571 37703 28577
rect 37734 28568 37740 28580
rect 37792 28568 37798 28620
rect 18509 28543 18567 28549
rect 18509 28509 18521 28543
rect 18555 28509 18567 28543
rect 18509 28503 18567 28509
rect 20349 28543 20407 28549
rect 20349 28509 20361 28543
rect 20395 28509 20407 28543
rect 20806 28540 20812 28552
rect 20767 28512 20812 28540
rect 20349 28503 20407 28509
rect 20806 28500 20812 28512
rect 20864 28500 20870 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 20990 28540 20996 28552
rect 20947 28512 20996 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 20990 28500 20996 28512
rect 21048 28500 21054 28552
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28509 21143 28543
rect 21085 28503 21143 28509
rect 11992 28472 12020 28500
rect 12161 28475 12219 28481
rect 12161 28472 12173 28475
rect 11992 28444 12173 28472
rect 12161 28441 12173 28444
rect 12207 28441 12219 28475
rect 12161 28435 12219 28441
rect 18693 28475 18751 28481
rect 18693 28441 18705 28475
rect 18739 28472 18751 28475
rect 19150 28472 19156 28484
rect 18739 28444 19156 28472
rect 18739 28441 18751 28444
rect 18693 28435 18751 28441
rect 19150 28432 19156 28444
rect 19208 28432 19214 28484
rect 20073 28475 20131 28481
rect 20073 28441 20085 28475
rect 20119 28472 20131 28475
rect 20162 28472 20168 28484
rect 20119 28444 20168 28472
rect 20119 28441 20131 28444
rect 20073 28435 20131 28441
rect 20162 28432 20168 28444
rect 20220 28432 20226 28484
rect 8573 28407 8631 28413
rect 8573 28373 8585 28407
rect 8619 28404 8631 28407
rect 8754 28404 8760 28416
rect 8619 28376 8760 28404
rect 8619 28373 8631 28376
rect 8573 28367 8631 28373
rect 8754 28364 8760 28376
rect 8812 28364 8818 28416
rect 11974 28413 11980 28416
rect 11961 28407 11980 28413
rect 11961 28373 11973 28407
rect 11961 28367 11980 28373
rect 11974 28364 11980 28367
rect 12032 28364 12038 28416
rect 20257 28407 20315 28413
rect 20257 28373 20269 28407
rect 20303 28404 20315 28407
rect 20898 28404 20904 28416
rect 20303 28376 20904 28404
rect 20303 28373 20315 28376
rect 20257 28367 20315 28373
rect 20898 28364 20904 28376
rect 20956 28364 20962 28416
rect 21100 28404 21128 28503
rect 21174 28500 21180 28552
rect 21232 28540 21238 28552
rect 21818 28540 21824 28552
rect 21232 28512 21277 28540
rect 21779 28512 21824 28540
rect 21232 28500 21238 28512
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 25222 28540 25228 28552
rect 25183 28512 25228 28540
rect 25222 28500 25228 28512
rect 25280 28500 25286 28552
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28540 28043 28543
rect 28534 28540 28540 28552
rect 28031 28512 28540 28540
rect 28031 28509 28043 28512
rect 27985 28503 28043 28509
rect 28534 28500 28540 28512
rect 28592 28500 28598 28552
rect 28994 28500 29000 28552
rect 29052 28540 29058 28552
rect 29825 28543 29883 28549
rect 29825 28540 29837 28543
rect 29052 28512 29837 28540
rect 29052 28500 29058 28512
rect 29825 28509 29837 28512
rect 29871 28540 29883 28543
rect 30190 28540 30196 28552
rect 29871 28512 30196 28540
rect 29871 28509 29883 28512
rect 29825 28503 29883 28509
rect 30190 28500 30196 28512
rect 30248 28500 30254 28552
rect 31386 28500 31392 28552
rect 31444 28540 31450 28552
rect 31665 28543 31723 28549
rect 31665 28540 31677 28543
rect 31444 28512 31677 28540
rect 31444 28500 31450 28512
rect 31665 28509 31677 28512
rect 31711 28509 31723 28543
rect 31665 28503 31723 28509
rect 35250 28500 35256 28552
rect 35308 28540 35314 28552
rect 35805 28543 35863 28549
rect 35805 28540 35817 28543
rect 35308 28512 35817 28540
rect 35308 28500 35314 28512
rect 35805 28509 35817 28512
rect 35851 28509 35863 28543
rect 35805 28503 35863 28509
rect 37918 28500 37924 28552
rect 37976 28540 37982 28552
rect 38105 28543 38163 28549
rect 38105 28540 38117 28543
rect 37976 28512 38117 28540
rect 37976 28500 37982 28512
rect 38105 28509 38117 28512
rect 38151 28509 38163 28543
rect 38105 28503 38163 28509
rect 25498 28481 25504 28484
rect 21361 28475 21419 28481
rect 21361 28441 21373 28475
rect 21407 28472 21419 28475
rect 22066 28475 22124 28481
rect 22066 28472 22078 28475
rect 21407 28444 22078 28472
rect 21407 28441 21419 28444
rect 21361 28435 21419 28441
rect 22066 28441 22078 28444
rect 22112 28441 22124 28475
rect 22066 28435 22124 28441
rect 23032 28444 25452 28472
rect 23032 28404 23060 28444
rect 23198 28404 23204 28416
rect 21100 28376 23060 28404
rect 23111 28376 23204 28404
rect 23198 28364 23204 28376
rect 23256 28404 23262 28416
rect 24394 28404 24400 28416
rect 23256 28376 24400 28404
rect 23256 28364 23262 28376
rect 24394 28364 24400 28376
rect 24452 28364 24458 28416
rect 25424 28404 25452 28444
rect 25492 28435 25504 28481
rect 25556 28472 25562 28484
rect 25556 28444 25592 28472
rect 25498 28432 25504 28435
rect 25556 28432 25562 28444
rect 30374 28432 30380 28484
rect 30432 28472 30438 28484
rect 31021 28475 31079 28481
rect 31021 28472 31033 28475
rect 30432 28444 31033 28472
rect 30432 28432 30438 28444
rect 31021 28441 31033 28444
rect 31067 28472 31079 28475
rect 31757 28475 31815 28481
rect 31757 28472 31769 28475
rect 31067 28444 31769 28472
rect 31067 28441 31079 28444
rect 31021 28435 31079 28441
rect 31757 28441 31769 28444
rect 31803 28441 31815 28475
rect 35986 28472 35992 28484
rect 35947 28444 35992 28472
rect 31757 28435 31815 28441
rect 35986 28432 35992 28444
rect 36044 28432 36050 28484
rect 37734 28432 37740 28484
rect 37792 28472 37798 28484
rect 38194 28472 38200 28484
rect 37792 28444 38200 28472
rect 37792 28432 37798 28444
rect 38194 28432 38200 28444
rect 38252 28432 38258 28484
rect 26326 28404 26332 28416
rect 25424 28376 26332 28404
rect 26326 28364 26332 28376
rect 26384 28364 26390 28416
rect 27798 28404 27804 28416
rect 27759 28376 27804 28404
rect 27798 28364 27804 28376
rect 27856 28364 27862 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 12253 28203 12311 28209
rect 12253 28169 12265 28203
rect 12299 28169 12311 28203
rect 12253 28163 12311 28169
rect 15197 28203 15255 28209
rect 15197 28169 15209 28203
rect 15243 28200 15255 28203
rect 19886 28200 19892 28212
rect 15243 28172 17264 28200
rect 15243 28169 15255 28172
rect 15197 28163 15255 28169
rect 12268 28132 12296 28163
rect 12268 28104 16068 28132
rect 1854 28064 1860 28076
rect 1815 28036 1860 28064
rect 1854 28024 1860 28036
rect 1912 28024 1918 28076
rect 4246 28024 4252 28076
rect 4304 28064 4310 28076
rect 4341 28067 4399 28073
rect 4341 28064 4353 28067
rect 4304 28036 4353 28064
rect 4304 28024 4310 28036
rect 4341 28033 4353 28036
rect 4387 28033 4399 28067
rect 8846 28064 8852 28076
rect 8807 28036 8852 28064
rect 4341 28027 4399 28033
rect 8846 28024 8852 28036
rect 8904 28024 8910 28076
rect 11146 28024 11152 28076
rect 11204 28064 11210 28076
rect 11885 28067 11943 28073
rect 11885 28064 11897 28067
rect 11204 28036 11897 28064
rect 11204 28024 11210 28036
rect 11885 28033 11897 28036
rect 11931 28033 11943 28067
rect 13262 28064 13268 28076
rect 13223 28036 13268 28064
rect 11885 28027 11943 28033
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 14752 28073 14780 28104
rect 14737 28067 14795 28073
rect 14737 28033 14749 28067
rect 14783 28033 14795 28067
rect 15197 28067 15255 28073
rect 15197 28064 15209 28067
rect 14737 28027 14795 28033
rect 14844 28036 15209 28064
rect 2038 27996 2044 28008
rect 1999 27968 2044 27996
rect 2038 27956 2044 27968
rect 2096 27956 2102 28008
rect 2774 27996 2780 28008
rect 2735 27968 2780 27996
rect 2774 27956 2780 27968
rect 2832 27956 2838 28008
rect 8754 27996 8760 28008
rect 8715 27968 8760 27996
rect 8754 27956 8760 27968
rect 8812 27956 8818 28008
rect 11790 27996 11796 28008
rect 11751 27968 11796 27996
rect 11790 27956 11796 27968
rect 11848 27956 11854 28008
rect 13354 27996 13360 28008
rect 13315 27968 13360 27996
rect 13354 27956 13360 27968
rect 13412 27956 13418 28008
rect 14844 27996 14872 28036
rect 15197 28033 15209 28036
rect 15243 28064 15255 28067
rect 15378 28064 15384 28076
rect 15243 28036 15384 28064
rect 15243 28033 15255 28036
rect 15197 28027 15255 28033
rect 15378 28024 15384 28036
rect 15436 28064 15442 28076
rect 16040 28073 16068 28104
rect 16206 28092 16212 28144
rect 16264 28132 16270 28144
rect 17236 28141 17264 28172
rect 19306 28172 19892 28200
rect 17005 28135 17063 28141
rect 17005 28132 17017 28135
rect 16264 28104 17017 28132
rect 16264 28092 16270 28104
rect 17005 28101 17017 28104
rect 17051 28101 17063 28135
rect 17005 28095 17063 28101
rect 17221 28135 17279 28141
rect 17221 28101 17233 28135
rect 17267 28101 17279 28135
rect 17221 28095 17279 28101
rect 15933 28067 15991 28073
rect 15933 28064 15945 28067
rect 15436 28036 15945 28064
rect 15436 28024 15442 28036
rect 15933 28033 15945 28036
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 16025 28067 16083 28073
rect 16025 28033 16037 28067
rect 16071 28033 16083 28067
rect 16025 28027 16083 28033
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28033 16175 28067
rect 16117 28027 16175 28033
rect 16301 28067 16359 28073
rect 16301 28033 16313 28067
rect 16347 28064 16359 28067
rect 19306 28064 19334 28172
rect 19886 28160 19892 28172
rect 19944 28200 19950 28212
rect 22922 28200 22928 28212
rect 19944 28172 22928 28200
rect 19944 28160 19950 28172
rect 22922 28160 22928 28172
rect 22980 28160 22986 28212
rect 23553 28203 23611 28209
rect 23553 28169 23565 28203
rect 23599 28200 23611 28203
rect 24026 28200 24032 28212
rect 23599 28172 24032 28200
rect 23599 28169 23611 28172
rect 23553 28163 23611 28169
rect 24026 28160 24032 28172
rect 24084 28160 24090 28212
rect 26418 28200 26424 28212
rect 25976 28172 26424 28200
rect 20254 28132 20260 28144
rect 16347 28036 19334 28064
rect 19628 28104 20260 28132
rect 16347 28033 16359 28036
rect 16301 28027 16359 28033
rect 14752 27968 14872 27996
rect 15013 27999 15071 28005
rect 11054 27888 11060 27940
rect 11112 27928 11118 27940
rect 12897 27931 12955 27937
rect 12897 27928 12909 27931
rect 11112 27900 12909 27928
rect 11112 27888 11118 27900
rect 12897 27897 12909 27900
rect 12943 27897 12955 27931
rect 12897 27891 12955 27897
rect 9125 27863 9183 27869
rect 9125 27829 9137 27863
rect 9171 27860 9183 27863
rect 14752 27860 14780 27968
rect 15013 27965 15025 27999
rect 15059 27996 15071 27999
rect 15562 27996 15568 28008
rect 15059 27968 15568 27996
rect 15059 27965 15071 27968
rect 15013 27959 15071 27965
rect 15562 27956 15568 27968
rect 15620 27956 15626 28008
rect 16132 27996 16160 28027
rect 19628 27996 19656 28104
rect 20254 28092 20260 28104
rect 20312 28132 20318 28144
rect 20533 28135 20591 28141
rect 20533 28132 20545 28135
rect 20312 28104 20545 28132
rect 20312 28092 20318 28104
rect 20533 28101 20545 28104
rect 20579 28101 20591 28135
rect 23750 28132 23756 28144
rect 20533 28095 20591 28101
rect 22756 28104 23336 28132
rect 23711 28104 23756 28132
rect 22756 28076 22784 28104
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 19981 28067 20039 28073
rect 19981 28033 19993 28067
rect 20027 28064 20039 28067
rect 20162 28064 20168 28076
rect 20027 28036 20168 28064
rect 20027 28033 20039 28036
rect 19981 28027 20039 28033
rect 16132 27968 19656 27996
rect 15657 27931 15715 27937
rect 15657 27897 15669 27931
rect 15703 27928 15715 27931
rect 15703 27900 17080 27928
rect 15703 27897 15715 27900
rect 15657 27891 15715 27897
rect 9171 27832 14780 27860
rect 14875 27863 14933 27869
rect 9171 27829 9183 27832
rect 9125 27823 9183 27829
rect 14875 27829 14887 27863
rect 14921 27860 14933 27863
rect 15746 27860 15752 27872
rect 14921 27832 15752 27860
rect 14921 27829 14933 27832
rect 14875 27823 14933 27829
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 16850 27860 16856 27872
rect 16811 27832 16856 27860
rect 16850 27820 16856 27832
rect 16908 27820 16914 27872
rect 17052 27869 17080 27900
rect 17678 27888 17684 27940
rect 17736 27928 17742 27940
rect 19720 27928 19748 28027
rect 20162 28024 20168 28036
rect 20220 28024 20226 28076
rect 22738 28064 22744 28076
rect 22699 28036 22744 28064
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 22925 28067 22983 28073
rect 22925 28033 22937 28067
rect 22971 28064 22983 28067
rect 23198 28064 23204 28076
rect 22971 28036 23204 28064
rect 22971 28033 22983 28036
rect 22925 28027 22983 28033
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23308 28064 23336 28104
rect 23750 28092 23756 28104
rect 23808 28092 23814 28144
rect 24581 28135 24639 28141
rect 24581 28132 24593 28135
rect 23860 28104 24593 28132
rect 23860 28064 23888 28104
rect 24581 28101 24593 28104
rect 24627 28101 24639 28135
rect 24581 28095 24639 28101
rect 24394 28064 24400 28076
rect 23308 28036 23888 28064
rect 24307 28036 24400 28064
rect 24394 28024 24400 28036
rect 24452 28064 24458 28076
rect 25976 28064 26004 28172
rect 26418 28160 26424 28172
rect 26476 28160 26482 28212
rect 29086 28160 29092 28212
rect 29144 28200 29150 28212
rect 29273 28203 29331 28209
rect 29273 28200 29285 28203
rect 29144 28172 29285 28200
rect 29144 28160 29150 28172
rect 29273 28169 29285 28172
rect 29319 28169 29331 28203
rect 32306 28200 32312 28212
rect 29273 28163 29331 28169
rect 29380 28172 31754 28200
rect 32267 28172 32312 28200
rect 29380 28132 29408 28172
rect 24452 28036 26004 28064
rect 26068 28104 29408 28132
rect 30377 28135 30435 28141
rect 24452 28024 24458 28036
rect 19889 27999 19947 28005
rect 19889 27965 19901 27999
rect 19935 27996 19947 27999
rect 20070 27996 20076 28008
rect 19935 27968 20076 27996
rect 19935 27965 19947 27968
rect 19889 27959 19947 27965
rect 20070 27956 20076 27968
rect 20128 27956 20134 28008
rect 20993 27999 21051 28005
rect 20993 27965 21005 27999
rect 21039 27996 21051 27999
rect 26068 27996 26096 28104
rect 30377 28101 30389 28135
rect 30423 28132 30435 28135
rect 31726 28132 31754 28172
rect 32306 28160 32312 28172
rect 32364 28160 32370 28212
rect 35250 28200 35256 28212
rect 35211 28172 35256 28200
rect 35250 28160 35256 28172
rect 35308 28160 35314 28212
rect 35986 28200 35992 28212
rect 35947 28172 35992 28200
rect 35986 28160 35992 28172
rect 36044 28160 36050 28212
rect 30423 28104 30972 28132
rect 31726 28104 35112 28132
rect 30423 28101 30435 28104
rect 30377 28095 30435 28101
rect 26145 28067 26203 28073
rect 26145 28033 26157 28067
rect 26191 28064 26203 28067
rect 26326 28064 26332 28076
rect 26191 28036 26332 28064
rect 26191 28033 26203 28036
rect 26145 28027 26203 28033
rect 26326 28024 26332 28036
rect 26384 28064 26390 28076
rect 26970 28064 26976 28076
rect 26384 28036 26976 28064
rect 26384 28024 26390 28036
rect 26970 28024 26976 28036
rect 27028 28024 27034 28076
rect 28166 28073 28172 28076
rect 28160 28027 28172 28073
rect 28224 28064 28230 28076
rect 30101 28067 30159 28073
rect 28224 28036 28260 28064
rect 28166 28024 28172 28027
rect 28224 28024 28230 28036
rect 30101 28033 30113 28067
rect 30147 28033 30159 28067
rect 30101 28027 30159 28033
rect 21039 27968 26096 27996
rect 26237 27999 26295 28005
rect 21039 27965 21051 27968
rect 20993 27959 21051 27965
rect 26237 27965 26249 27999
rect 26283 27996 26295 27999
rect 26510 27996 26516 28008
rect 26283 27968 26516 27996
rect 26283 27965 26295 27968
rect 26237 27959 26295 27965
rect 26510 27956 26516 27968
rect 26568 27956 26574 28008
rect 27893 27999 27951 28005
rect 27893 27965 27905 27999
rect 27939 27965 27951 27999
rect 27893 27959 27951 27965
rect 17736 27900 19748 27928
rect 19797 27931 19855 27937
rect 17736 27888 17742 27900
rect 19797 27897 19809 27931
rect 19843 27928 19855 27931
rect 19978 27928 19984 27940
rect 19843 27900 19984 27928
rect 19843 27897 19855 27900
rect 19797 27891 19855 27897
rect 19978 27888 19984 27900
rect 20036 27888 20042 27940
rect 20254 27888 20260 27940
rect 20312 27928 20318 27940
rect 20809 27931 20867 27937
rect 20809 27928 20821 27931
rect 20312 27900 20821 27928
rect 20312 27888 20318 27900
rect 20809 27897 20821 27900
rect 20855 27897 20867 27931
rect 20809 27891 20867 27897
rect 23032 27900 23612 27928
rect 23032 27872 23060 27900
rect 17037 27863 17095 27869
rect 17037 27829 17049 27863
rect 17083 27829 17095 27863
rect 17037 27823 17095 27829
rect 19521 27863 19579 27869
rect 19521 27829 19533 27863
rect 19567 27860 19579 27863
rect 19610 27860 19616 27872
rect 19567 27832 19616 27860
rect 19567 27829 19579 27832
rect 19521 27823 19579 27829
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 22833 27863 22891 27869
rect 22833 27829 22845 27863
rect 22879 27860 22891 27863
rect 23014 27860 23020 27872
rect 22879 27832 23020 27860
rect 22879 27829 22891 27832
rect 22833 27823 22891 27829
rect 23014 27820 23020 27832
rect 23072 27820 23078 27872
rect 23385 27863 23443 27869
rect 23385 27829 23397 27863
rect 23431 27860 23443 27863
rect 23474 27860 23480 27872
rect 23431 27832 23480 27860
rect 23431 27829 23443 27832
rect 23385 27823 23443 27829
rect 23474 27820 23480 27832
rect 23532 27820 23538 27872
rect 23584 27869 23612 27900
rect 25222 27888 25228 27940
rect 25280 27928 25286 27940
rect 27908 27928 27936 27959
rect 25280 27900 27936 27928
rect 30116 27928 30144 28027
rect 30190 28024 30196 28076
rect 30248 28064 30254 28076
rect 30944 28073 30972 28104
rect 30929 28067 30987 28073
rect 30248 28036 30293 28064
rect 30248 28024 30254 28036
rect 30929 28033 30941 28067
rect 30975 28033 30987 28067
rect 30929 28027 30987 28033
rect 31018 28024 31024 28076
rect 31076 28064 31082 28076
rect 31205 28067 31263 28073
rect 31076 28036 31121 28064
rect 31076 28024 31082 28036
rect 31205 28033 31217 28067
rect 31251 28064 31263 28067
rect 31754 28064 31760 28076
rect 31251 28036 31760 28064
rect 31251 28033 31263 28036
rect 31205 28027 31263 28033
rect 31754 28024 31760 28036
rect 31812 28024 31818 28076
rect 35084 28073 35112 28104
rect 32493 28067 32551 28073
rect 32493 28033 32505 28067
rect 32539 28033 32551 28067
rect 32493 28027 32551 28033
rect 35069 28067 35127 28073
rect 35069 28033 35081 28067
rect 35115 28033 35127 28067
rect 35069 28027 35127 28033
rect 35897 28067 35955 28073
rect 35897 28033 35909 28067
rect 35943 28064 35955 28067
rect 36446 28064 36452 28076
rect 35943 28036 36452 28064
rect 35943 28033 35955 28036
rect 35897 28027 35955 28033
rect 30374 27996 30380 28008
rect 30335 27968 30380 27996
rect 30374 27956 30380 27968
rect 30432 27956 30438 28008
rect 31113 27999 31171 28005
rect 31113 27965 31125 27999
rect 31159 27996 31171 27999
rect 31662 27996 31668 28008
rect 31159 27968 31668 27996
rect 31159 27965 31171 27968
rect 31113 27959 31171 27965
rect 31662 27956 31668 27968
rect 31720 27996 31726 28008
rect 32508 27996 32536 28027
rect 36446 28024 36452 28036
rect 36504 28024 36510 28076
rect 31720 27968 32536 27996
rect 32677 27999 32735 28005
rect 31720 27956 31726 27968
rect 32677 27965 32689 27999
rect 32723 27965 32735 27999
rect 32677 27959 32735 27965
rect 30116 27900 31156 27928
rect 25280 27888 25286 27900
rect 31128 27872 31156 27900
rect 31754 27888 31760 27940
rect 31812 27928 31818 27940
rect 32692 27928 32720 27959
rect 31812 27900 32720 27928
rect 31812 27888 31818 27900
rect 23569 27863 23627 27869
rect 23569 27829 23581 27863
rect 23615 27829 23627 27863
rect 23569 27823 23627 27829
rect 24026 27820 24032 27872
rect 24084 27860 24090 27872
rect 24213 27863 24271 27869
rect 24213 27860 24225 27863
rect 24084 27832 24225 27860
rect 24084 27820 24090 27832
rect 24213 27829 24225 27832
rect 24259 27829 24271 27863
rect 24213 27823 24271 27829
rect 25777 27863 25835 27869
rect 25777 27829 25789 27863
rect 25823 27860 25835 27863
rect 26234 27860 26240 27872
rect 25823 27832 26240 27860
rect 25823 27829 25835 27832
rect 25777 27823 25835 27829
rect 26234 27820 26240 27832
rect 26292 27820 26298 27872
rect 31110 27820 31116 27872
rect 31168 27820 31174 27872
rect 31389 27863 31447 27869
rect 31389 27829 31401 27863
rect 31435 27860 31447 27863
rect 31478 27860 31484 27872
rect 31435 27832 31484 27860
rect 31435 27829 31447 27832
rect 31389 27823 31447 27829
rect 31478 27820 31484 27832
rect 31536 27820 31542 27872
rect 36446 27820 36452 27872
rect 36504 27860 36510 27872
rect 37553 27863 37611 27869
rect 37553 27860 37565 27863
rect 36504 27832 37565 27860
rect 36504 27820 36510 27832
rect 37553 27829 37565 27832
rect 37599 27829 37611 27863
rect 37553 27823 37611 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2038 27616 2044 27668
rect 2096 27656 2102 27668
rect 2133 27659 2191 27665
rect 2133 27656 2145 27659
rect 2096 27628 2145 27656
rect 2096 27616 2102 27628
rect 2133 27625 2145 27628
rect 2179 27625 2191 27659
rect 11790 27656 11796 27668
rect 2133 27619 2191 27625
rect 10980 27628 11796 27656
rect 9861 27591 9919 27597
rect 9861 27557 9873 27591
rect 9907 27588 9919 27591
rect 10980 27588 11008 27628
rect 11790 27616 11796 27628
rect 11848 27616 11854 27668
rect 15933 27659 15991 27665
rect 15933 27625 15945 27659
rect 15979 27656 15991 27659
rect 16206 27656 16212 27668
rect 15979 27628 16212 27656
rect 15979 27625 15991 27628
rect 15933 27619 15991 27625
rect 16206 27616 16212 27628
rect 16264 27616 16270 27668
rect 19886 27656 19892 27668
rect 19847 27628 19892 27656
rect 19886 27616 19892 27628
rect 19944 27616 19950 27668
rect 20993 27659 21051 27665
rect 20993 27625 21005 27659
rect 21039 27625 21051 27659
rect 20993 27619 21051 27625
rect 30561 27659 30619 27665
rect 30561 27625 30573 27659
rect 30607 27656 30619 27659
rect 31018 27656 31024 27668
rect 30607 27628 31024 27656
rect 30607 27625 30619 27628
rect 30561 27619 30619 27625
rect 11146 27588 11152 27600
rect 9907 27560 11008 27588
rect 11107 27560 11152 27588
rect 9907 27557 9919 27560
rect 9861 27551 9919 27557
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 13354 27588 13360 27600
rect 13315 27560 13360 27588
rect 13354 27548 13360 27560
rect 13412 27548 13418 27600
rect 9582 27520 9588 27532
rect 9543 27492 9588 27520
rect 9582 27480 9588 27492
rect 9640 27480 9646 27532
rect 10873 27523 10931 27529
rect 10873 27489 10885 27523
rect 10919 27520 10931 27523
rect 11054 27520 11060 27532
rect 10919 27492 11060 27520
rect 10919 27489 10931 27492
rect 10873 27483 10931 27489
rect 11054 27480 11060 27492
rect 11112 27480 11118 27532
rect 13078 27520 13084 27532
rect 13039 27492 13084 27520
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 18414 27520 18420 27532
rect 18375 27492 18420 27520
rect 18414 27480 18420 27492
rect 18472 27480 18478 27532
rect 19426 27520 19432 27532
rect 19387 27492 19432 27520
rect 19426 27480 19432 27492
rect 19484 27480 19490 27532
rect 21008 27520 21036 27619
rect 31018 27616 31024 27628
rect 31076 27616 31082 27668
rect 31662 27616 31668 27668
rect 31720 27656 31726 27668
rect 31757 27659 31815 27665
rect 31757 27656 31769 27659
rect 31720 27628 31769 27656
rect 31720 27616 31726 27628
rect 31757 27625 31769 27628
rect 31803 27625 31815 27659
rect 31757 27619 31815 27625
rect 27525 27591 27583 27597
rect 27525 27557 27537 27591
rect 27571 27588 27583 27591
rect 27798 27588 27804 27600
rect 27571 27560 27804 27588
rect 27571 27557 27583 27560
rect 27525 27551 27583 27557
rect 27798 27548 27804 27560
rect 27856 27548 27862 27600
rect 27982 27548 27988 27600
rect 28040 27588 28046 27600
rect 28534 27588 28540 27600
rect 28040 27560 28540 27588
rect 28040 27548 28046 27560
rect 28534 27548 28540 27560
rect 28592 27548 28598 27600
rect 21266 27520 21272 27532
rect 21008 27492 21272 27520
rect 21266 27480 21272 27492
rect 21324 27480 21330 27532
rect 23569 27523 23627 27529
rect 23569 27520 23581 27523
rect 23032 27492 23581 27520
rect 23032 27464 23060 27492
rect 23569 27489 23581 27492
rect 23615 27489 23627 27523
rect 27430 27520 27436 27532
rect 23569 27483 23627 27489
rect 26712 27492 27436 27520
rect 26712 27464 26740 27492
rect 27430 27480 27436 27492
rect 27488 27480 27494 27532
rect 30374 27480 30380 27532
rect 30432 27520 30438 27532
rect 30432 27492 30788 27520
rect 30432 27480 30438 27492
rect 2225 27455 2283 27461
rect 2225 27421 2237 27455
rect 2271 27452 2283 27455
rect 2406 27452 2412 27464
rect 2271 27424 2412 27452
rect 2271 27421 2283 27424
rect 2225 27415 2283 27421
rect 2406 27412 2412 27424
rect 2464 27452 2470 27464
rect 3602 27452 3608 27464
rect 2464 27424 3608 27452
rect 2464 27412 2470 27424
rect 3602 27412 3608 27424
rect 3660 27412 3666 27464
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 9493 27455 9551 27461
rect 9493 27452 9505 27455
rect 9456 27424 9505 27452
rect 9456 27412 9462 27424
rect 9493 27421 9505 27424
rect 9539 27421 9551 27455
rect 10778 27452 10784 27464
rect 10739 27424 10784 27452
rect 9493 27415 9551 27421
rect 10778 27412 10784 27424
rect 10836 27412 10842 27464
rect 12989 27455 13047 27461
rect 12989 27421 13001 27455
rect 13035 27452 13047 27455
rect 13906 27452 13912 27464
rect 13035 27424 13912 27452
rect 13035 27421 13047 27424
rect 12989 27415 13047 27421
rect 13906 27412 13912 27424
rect 13964 27412 13970 27464
rect 15378 27452 15384 27464
rect 15339 27424 15384 27452
rect 15378 27412 15384 27424
rect 15436 27412 15442 27464
rect 15470 27412 15476 27464
rect 15528 27452 15534 27464
rect 15654 27452 15660 27464
rect 15528 27424 15573 27452
rect 15615 27424 15660 27452
rect 15528 27412 15534 27424
rect 15654 27412 15660 27424
rect 15712 27412 15718 27464
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 19610 27452 19616 27464
rect 15804 27424 15849 27452
rect 19571 27424 19616 27452
rect 15804 27412 15810 27424
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 19981 27455 20039 27461
rect 19981 27421 19993 27455
rect 20027 27452 20039 27455
rect 20254 27452 20260 27464
rect 20027 27424 20260 27452
rect 20027 27421 20039 27424
rect 19981 27415 20039 27421
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 20990 27412 20996 27464
rect 21048 27452 21054 27464
rect 23014 27452 23020 27464
rect 21048 27424 21220 27452
rect 22975 27424 23020 27452
rect 21048 27412 21054 27424
rect 18138 27384 18144 27396
rect 18196 27393 18202 27396
rect 18108 27356 18144 27384
rect 18138 27344 18144 27356
rect 18196 27347 18208 27393
rect 20809 27387 20867 27393
rect 20809 27353 20821 27387
rect 20855 27384 20867 27387
rect 20898 27384 20904 27396
rect 20855 27356 20904 27384
rect 20855 27353 20867 27356
rect 20809 27347 20867 27353
rect 18196 27344 18202 27347
rect 20898 27344 20904 27356
rect 20956 27344 20962 27396
rect 15654 27276 15660 27328
rect 15712 27316 15718 27328
rect 17037 27319 17095 27325
rect 17037 27316 17049 27319
rect 15712 27288 17049 27316
rect 15712 27276 15718 27288
rect 17037 27285 17049 27288
rect 17083 27285 17095 27319
rect 17037 27279 17095 27285
rect 19426 27276 19432 27328
rect 19484 27316 19490 27328
rect 21192 27325 21220 27424
rect 23014 27412 23020 27424
rect 23072 27412 23078 27464
rect 23109 27455 23167 27461
rect 23109 27421 23121 27455
rect 23155 27452 23167 27455
rect 24026 27452 24032 27464
rect 23155 27424 24032 27452
rect 23155 27421 23167 27424
rect 23109 27415 23167 27421
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27421 25191 27455
rect 25133 27415 25191 27421
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27452 25375 27455
rect 26694 27452 26700 27464
rect 25363 27424 26700 27452
rect 25363 27421 25375 27424
rect 25317 27415 25375 27421
rect 22833 27387 22891 27393
rect 22833 27353 22845 27387
rect 22879 27384 22891 27387
rect 23566 27384 23572 27396
rect 22879 27356 23572 27384
rect 22879 27353 22891 27356
rect 22833 27347 22891 27353
rect 23566 27344 23572 27356
rect 23624 27384 23630 27396
rect 23750 27384 23756 27396
rect 23624 27356 23756 27384
rect 23624 27344 23630 27356
rect 23750 27344 23756 27356
rect 23808 27344 23814 27396
rect 24854 27344 24860 27396
rect 24912 27384 24918 27396
rect 25148 27384 25176 27415
rect 26694 27412 26700 27424
rect 26752 27412 26758 27464
rect 27338 27452 27344 27464
rect 27251 27424 27344 27452
rect 27338 27412 27344 27424
rect 27396 27452 27402 27464
rect 27522 27452 27528 27464
rect 27396 27424 27528 27452
rect 27396 27412 27402 27424
rect 27522 27412 27528 27424
rect 27580 27412 27586 27464
rect 27617 27455 27675 27461
rect 27617 27421 27629 27455
rect 27663 27452 27675 27455
rect 27706 27452 27712 27464
rect 27663 27424 27712 27452
rect 27663 27421 27675 27424
rect 27617 27415 27675 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 28721 27455 28779 27461
rect 28721 27421 28733 27455
rect 28767 27452 28779 27455
rect 29086 27452 29092 27464
rect 28767 27424 29092 27452
rect 28767 27421 28779 27424
rect 28721 27415 28779 27421
rect 29086 27412 29092 27424
rect 29144 27412 29150 27464
rect 30190 27412 30196 27464
rect 30248 27452 30254 27464
rect 30760 27461 30788 27492
rect 31110 27480 31116 27532
rect 31168 27520 31174 27532
rect 31297 27523 31355 27529
rect 31297 27520 31309 27523
rect 31168 27492 31309 27520
rect 31168 27480 31174 27492
rect 31297 27489 31309 27492
rect 31343 27489 31355 27523
rect 31297 27483 31355 27489
rect 30561 27455 30619 27461
rect 30561 27452 30573 27455
rect 30248 27424 30573 27452
rect 30248 27412 30254 27424
rect 30561 27421 30573 27424
rect 30607 27421 30619 27455
rect 30561 27415 30619 27421
rect 30745 27455 30803 27461
rect 30745 27421 30757 27455
rect 30791 27421 30803 27455
rect 31386 27452 31392 27464
rect 31347 27424 31392 27452
rect 30745 27415 30803 27421
rect 31386 27412 31392 27424
rect 31444 27412 31450 27464
rect 31772 27452 31800 27619
rect 32309 27523 32367 27529
rect 32309 27489 32321 27523
rect 32355 27520 32367 27523
rect 32490 27520 32496 27532
rect 32355 27492 32496 27520
rect 32355 27489 32367 27492
rect 32309 27483 32367 27489
rect 32490 27480 32496 27492
rect 32548 27480 32554 27532
rect 36446 27520 36452 27532
rect 36407 27492 36452 27520
rect 36446 27480 36452 27492
rect 36504 27480 36510 27532
rect 32217 27455 32275 27461
rect 32217 27452 32229 27455
rect 31772 27424 32229 27452
rect 32217 27421 32229 27424
rect 32263 27421 32275 27455
rect 32217 27415 32275 27421
rect 32401 27455 32459 27461
rect 32401 27421 32413 27455
rect 32447 27421 32459 27455
rect 32401 27415 32459 27421
rect 26050 27384 26056 27396
rect 24912 27356 26056 27384
rect 24912 27344 24918 27356
rect 26050 27344 26056 27356
rect 26108 27384 26114 27396
rect 30650 27384 30656 27396
rect 26108 27356 30656 27384
rect 26108 27344 26114 27356
rect 30650 27344 30656 27356
rect 30708 27344 30714 27396
rect 31754 27344 31760 27396
rect 31812 27384 31818 27396
rect 32416 27384 32444 27415
rect 31812 27356 32444 27384
rect 36633 27387 36691 27393
rect 31812 27344 31818 27356
rect 36633 27353 36645 27387
rect 36679 27384 36691 27387
rect 37550 27384 37556 27396
rect 36679 27356 37556 27384
rect 36679 27353 36691 27356
rect 36633 27347 36691 27353
rect 37550 27344 37556 27356
rect 37608 27344 37614 27396
rect 38286 27384 38292 27396
rect 38247 27356 38292 27384
rect 38286 27344 38292 27356
rect 38344 27344 38350 27396
rect 21009 27319 21067 27325
rect 21009 27316 21021 27319
rect 19484 27288 21021 27316
rect 19484 27276 19490 27288
rect 21009 27285 21021 27288
rect 21055 27285 21067 27319
rect 21009 27279 21067 27285
rect 21177 27319 21235 27325
rect 21177 27285 21189 27319
rect 21223 27316 21235 27319
rect 21726 27316 21732 27328
rect 21223 27288 21732 27316
rect 21223 27285 21235 27288
rect 21177 27279 21235 27285
rect 21726 27276 21732 27288
rect 21784 27276 21790 27328
rect 22922 27276 22928 27328
rect 22980 27325 22986 27328
rect 22980 27316 22989 27325
rect 23842 27316 23848 27328
rect 22980 27288 23025 27316
rect 23803 27288 23848 27316
rect 22980 27279 22989 27288
rect 22980 27276 22986 27279
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 23937 27319 23995 27325
rect 23937 27285 23949 27319
rect 23983 27316 23995 27319
rect 24026 27316 24032 27328
rect 23983 27288 24032 27316
rect 23983 27285 23995 27288
rect 23937 27279 23995 27285
rect 24026 27276 24032 27288
rect 24084 27276 24090 27328
rect 25317 27319 25375 27325
rect 25317 27285 25329 27319
rect 25363 27316 25375 27319
rect 25682 27316 25688 27328
rect 25363 27288 25688 27316
rect 25363 27285 25375 27288
rect 25317 27279 25375 27285
rect 25682 27276 25688 27288
rect 25740 27276 25746 27328
rect 26418 27276 26424 27328
rect 26476 27316 26482 27328
rect 27157 27319 27215 27325
rect 27157 27316 27169 27319
rect 26476 27288 27169 27316
rect 26476 27276 26482 27288
rect 27157 27285 27169 27288
rect 27203 27285 27215 27319
rect 27157 27279 27215 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 18138 27072 18144 27124
rect 18196 27112 18202 27124
rect 18233 27115 18291 27121
rect 18233 27112 18245 27115
rect 18196 27084 18245 27112
rect 18196 27072 18202 27084
rect 18233 27081 18245 27084
rect 18279 27081 18291 27115
rect 18233 27075 18291 27081
rect 19061 27115 19119 27121
rect 19061 27081 19073 27115
rect 19107 27112 19119 27115
rect 20254 27112 20260 27124
rect 19107 27084 20260 27112
rect 19107 27081 19119 27084
rect 19061 27075 19119 27081
rect 20254 27072 20260 27084
rect 20312 27072 20318 27124
rect 25682 27112 25688 27124
rect 25643 27084 25688 27112
rect 25682 27072 25688 27084
rect 25740 27072 25746 27124
rect 37550 27112 37556 27124
rect 37511 27084 37556 27112
rect 37550 27072 37556 27084
rect 37608 27072 37614 27124
rect 16850 27044 16856 27056
rect 6886 27016 16856 27044
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 6886 26976 6914 27016
rect 16850 27004 16856 27016
rect 16908 27004 16914 27056
rect 17402 27044 17408 27056
rect 17363 27016 17408 27044
rect 17402 27004 17408 27016
rect 17460 27004 17466 27056
rect 22738 27004 22744 27056
rect 22796 27044 22802 27056
rect 22796 27016 23612 27044
rect 22796 27004 22802 27016
rect 8570 26976 8576 26988
rect 4295 26948 6914 26976
rect 8531 26948 8576 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 8757 26979 8815 26985
rect 8757 26945 8769 26979
rect 8803 26976 8815 26979
rect 8938 26976 8944 26988
rect 8803 26948 8944 26976
rect 8803 26945 8815 26948
rect 8757 26939 8815 26945
rect 8938 26936 8944 26948
rect 8996 26936 9002 26988
rect 9214 26976 9220 26988
rect 9175 26948 9220 26976
rect 9214 26936 9220 26948
rect 9272 26936 9278 26988
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26945 9459 26979
rect 9401 26939 9459 26945
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26976 11759 26979
rect 11885 26979 11943 26985
rect 11747 26948 11836 26976
rect 11747 26945 11759 26948
rect 11701 26939 11759 26945
rect 8665 26911 8723 26917
rect 8665 26877 8677 26911
rect 8711 26908 8723 26911
rect 9306 26908 9312 26920
rect 8711 26880 9312 26908
rect 8711 26877 8723 26880
rect 8665 26871 8723 26877
rect 9306 26868 9312 26880
rect 9364 26908 9370 26920
rect 9416 26908 9444 26939
rect 9364 26880 9444 26908
rect 9364 26868 9370 26880
rect 11808 26840 11836 26948
rect 11885 26945 11897 26979
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 11900 26908 11928 26939
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 12437 26979 12495 26985
rect 12437 26976 12449 26979
rect 12400 26948 12449 26976
rect 12400 26936 12406 26948
rect 12437 26945 12449 26948
rect 12483 26945 12495 26979
rect 12618 26976 12624 26988
rect 12579 26948 12624 26976
rect 12437 26939 12495 26945
rect 12618 26936 12624 26948
rect 12676 26936 12682 26988
rect 12802 26976 12808 26988
rect 12763 26948 12808 26976
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 18049 26979 18107 26985
rect 18049 26976 18061 26979
rect 17604 26948 18061 26976
rect 13906 26908 13912 26920
rect 11900 26880 13912 26908
rect 13906 26868 13912 26880
rect 13964 26868 13970 26920
rect 12710 26840 12716 26852
rect 11808 26812 12716 26840
rect 12710 26800 12716 26812
rect 12768 26800 12774 26852
rect 17037 26843 17095 26849
rect 17037 26840 17049 26843
rect 12820 26812 17049 26840
rect 3970 26732 3976 26784
rect 4028 26772 4034 26784
rect 4065 26775 4123 26781
rect 4065 26772 4077 26775
rect 4028 26744 4077 26772
rect 4028 26732 4034 26744
rect 4065 26741 4077 26744
rect 4111 26741 4123 26775
rect 9398 26772 9404 26784
rect 9359 26744 9404 26772
rect 4065 26735 4123 26741
rect 9398 26732 9404 26744
rect 9456 26732 9462 26784
rect 10870 26732 10876 26784
rect 10928 26772 10934 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 10928 26744 11805 26772
rect 10928 26732 10934 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 11793 26735 11851 26741
rect 11974 26732 11980 26784
rect 12032 26772 12038 26784
rect 12342 26772 12348 26784
rect 12032 26744 12348 26772
rect 12032 26732 12038 26744
rect 12342 26732 12348 26744
rect 12400 26772 12406 26784
rect 12820 26772 12848 26812
rect 17037 26809 17049 26812
rect 17083 26840 17095 26843
rect 17218 26840 17224 26852
rect 17083 26812 17224 26840
rect 17083 26809 17095 26812
rect 17037 26803 17095 26809
rect 17218 26800 17224 26812
rect 17276 26800 17282 26852
rect 17604 26849 17632 26948
rect 18049 26945 18061 26948
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 19061 26979 19119 26985
rect 19061 26945 19073 26979
rect 19107 26976 19119 26979
rect 19242 26976 19248 26988
rect 19107 26948 19248 26976
rect 19107 26945 19119 26948
rect 19061 26939 19119 26945
rect 19242 26936 19248 26948
rect 19300 26936 19306 26988
rect 23474 26976 23480 26988
rect 23435 26948 23480 26976
rect 23474 26936 23480 26948
rect 23532 26936 23538 26988
rect 23584 26976 23612 27016
rect 23842 27004 23848 27056
rect 23900 27044 23906 27056
rect 31754 27044 31760 27056
rect 23900 27016 31760 27044
rect 23900 27004 23906 27016
rect 31754 27004 31760 27016
rect 31812 27004 31818 27056
rect 24305 26979 24363 26985
rect 24305 26976 24317 26979
rect 23584 26948 24317 26976
rect 24305 26945 24317 26948
rect 24351 26945 24363 26979
rect 24305 26939 24363 26945
rect 24489 26979 24547 26985
rect 24489 26945 24501 26979
rect 24535 26976 24547 26979
rect 24854 26976 24860 26988
rect 24535 26948 24860 26976
rect 24535 26945 24547 26948
rect 24489 26939 24547 26945
rect 24854 26936 24860 26948
rect 24912 26936 24918 26988
rect 24946 26936 24952 26988
rect 25004 26976 25010 26988
rect 25501 26979 25559 26985
rect 25501 26976 25513 26979
rect 25004 26948 25513 26976
rect 25004 26936 25010 26948
rect 25501 26945 25513 26948
rect 25547 26945 25559 26979
rect 25501 26939 25559 26945
rect 25774 26936 25780 26988
rect 25832 26976 25838 26988
rect 26237 26979 26295 26985
rect 25832 26948 25877 26976
rect 25832 26936 25838 26948
rect 26237 26945 26249 26979
rect 26283 26945 26295 26979
rect 26237 26939 26295 26945
rect 26421 26979 26479 26985
rect 26421 26945 26433 26979
rect 26467 26976 26479 26979
rect 27338 26976 27344 26988
rect 26467 26948 27344 26976
rect 26467 26945 26479 26948
rect 26421 26939 26479 26945
rect 19334 26908 19340 26920
rect 19295 26880 19340 26908
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 23569 26911 23627 26917
rect 23569 26877 23581 26911
rect 23615 26908 23627 26911
rect 23934 26908 23940 26920
rect 23615 26880 23940 26908
rect 23615 26877 23627 26880
rect 23569 26871 23627 26877
rect 23934 26868 23940 26880
rect 23992 26868 23998 26920
rect 26252 26908 26280 26939
rect 27338 26936 27344 26948
rect 27396 26936 27402 26988
rect 27614 26936 27620 26988
rect 27672 26976 27678 26988
rect 27672 26948 29684 26976
rect 27672 26936 27678 26948
rect 27522 26908 27528 26920
rect 24872 26880 27528 26908
rect 24872 26852 24900 26880
rect 27522 26868 27528 26880
rect 27580 26868 27586 26920
rect 29270 26868 29276 26920
rect 29328 26908 29334 26920
rect 29549 26911 29607 26917
rect 29549 26908 29561 26911
rect 29328 26880 29561 26908
rect 29328 26868 29334 26880
rect 29549 26877 29561 26880
rect 29595 26877 29607 26911
rect 29656 26908 29684 26948
rect 29730 26936 29736 26988
rect 29788 26976 29794 26988
rect 29825 26979 29883 26985
rect 29825 26976 29837 26979
rect 29788 26948 29837 26976
rect 29788 26936 29794 26948
rect 29825 26945 29837 26948
rect 29871 26945 29883 26979
rect 37461 26979 37519 26985
rect 37461 26976 37473 26979
rect 29825 26939 29883 26945
rect 31726 26948 37473 26976
rect 31726 26908 31754 26948
rect 37461 26945 37473 26948
rect 37507 26945 37519 26979
rect 37461 26939 37519 26945
rect 29656 26880 31754 26908
rect 29549 26871 29607 26877
rect 17589 26843 17647 26849
rect 17589 26809 17601 26843
rect 17635 26809 17647 26843
rect 17589 26803 17647 26809
rect 18322 26800 18328 26852
rect 18380 26840 18386 26852
rect 19153 26843 19211 26849
rect 19153 26840 19165 26843
rect 18380 26812 19165 26840
rect 18380 26800 18386 26812
rect 19153 26809 19165 26812
rect 19199 26809 19211 26843
rect 19153 26803 19211 26809
rect 24854 26800 24860 26852
rect 24912 26800 24918 26852
rect 25498 26840 25504 26852
rect 25459 26812 25504 26840
rect 25498 26800 25504 26812
rect 25556 26800 25562 26852
rect 12400 26744 12848 26772
rect 12400 26732 12406 26744
rect 17310 26732 17316 26784
rect 17368 26772 17374 26784
rect 17405 26775 17463 26781
rect 17405 26772 17417 26775
rect 17368 26744 17417 26772
rect 17368 26732 17374 26744
rect 17405 26741 17417 26744
rect 17451 26772 17463 26775
rect 21358 26772 21364 26784
rect 17451 26744 21364 26772
rect 17451 26741 17463 26744
rect 17405 26735 17463 26741
rect 21358 26732 21364 26744
rect 21416 26732 21422 26784
rect 22922 26732 22928 26784
rect 22980 26772 22986 26784
rect 23477 26775 23535 26781
rect 23477 26772 23489 26775
rect 22980 26744 23489 26772
rect 22980 26732 22986 26744
rect 23477 26741 23489 26744
rect 23523 26741 23535 26775
rect 23477 26735 23535 26741
rect 23845 26775 23903 26781
rect 23845 26741 23857 26775
rect 23891 26772 23903 26775
rect 24302 26772 24308 26784
rect 23891 26744 24308 26772
rect 23891 26741 23903 26744
rect 23845 26735 23903 26741
rect 24302 26732 24308 26744
rect 24360 26732 24366 26784
rect 24397 26775 24455 26781
rect 24397 26741 24409 26775
rect 24443 26772 24455 26775
rect 24670 26772 24676 26784
rect 24443 26744 24676 26772
rect 24443 26741 24455 26744
rect 24397 26735 24455 26741
rect 24670 26732 24676 26744
rect 24728 26732 24734 26784
rect 26326 26772 26332 26784
rect 26287 26744 26332 26772
rect 26326 26732 26332 26744
rect 26384 26732 26390 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8754 26568 8760 26580
rect 8619 26540 8760 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 8754 26528 8760 26540
rect 8812 26568 8818 26580
rect 9214 26568 9220 26580
rect 8812 26540 9220 26568
rect 8812 26528 8818 26540
rect 9214 26528 9220 26540
rect 9272 26528 9278 26580
rect 9582 26568 9588 26580
rect 9543 26540 9588 26568
rect 9582 26528 9588 26540
rect 9640 26528 9646 26580
rect 10778 26528 10784 26580
rect 10836 26568 10842 26580
rect 12802 26568 12808 26580
rect 10836 26540 11192 26568
rect 12763 26540 12808 26568
rect 10836 26528 10842 26540
rect 4062 26460 4068 26512
rect 4120 26460 4126 26512
rect 11057 26503 11115 26509
rect 11057 26500 11069 26503
rect 9968 26472 11069 26500
rect 3970 26432 3976 26444
rect 3931 26404 3976 26432
rect 3970 26392 3976 26404
rect 4028 26392 4034 26444
rect 4080 26432 4108 26460
rect 4433 26435 4491 26441
rect 4433 26432 4445 26435
rect 4080 26404 4445 26432
rect 4433 26401 4445 26404
rect 4479 26401 4491 26435
rect 9398 26432 9404 26444
rect 9359 26404 9404 26432
rect 4433 26395 4491 26401
rect 9398 26392 9404 26404
rect 9456 26392 9462 26444
rect 8297 26367 8355 26373
rect 8297 26333 8309 26367
rect 8343 26333 8355 26367
rect 8297 26327 8355 26333
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 8938 26364 8944 26376
rect 8435 26336 8944 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 4154 26296 4160 26308
rect 4115 26268 4160 26296
rect 4154 26256 4160 26268
rect 4212 26256 4218 26308
rect 8312 26296 8340 26327
rect 8938 26324 8944 26336
rect 8996 26324 9002 26376
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26364 9367 26367
rect 9582 26364 9588 26376
rect 9355 26336 9588 26364
rect 9355 26333 9367 26336
rect 9309 26327 9367 26333
rect 9582 26324 9588 26336
rect 9640 26364 9646 26376
rect 9968 26364 9996 26472
rect 11057 26469 11069 26472
rect 11103 26469 11115 26503
rect 11057 26463 11115 26469
rect 11164 26432 11192 26540
rect 12802 26528 12808 26540
rect 12860 26528 12866 26580
rect 17402 26568 17408 26580
rect 17363 26540 17408 26568
rect 17402 26528 17408 26540
rect 17460 26528 17466 26580
rect 22557 26571 22615 26577
rect 22557 26537 22569 26571
rect 22603 26568 22615 26571
rect 22738 26568 22744 26580
rect 22603 26540 22744 26568
rect 22603 26537 22615 26540
rect 22557 26531 22615 26537
rect 22738 26528 22744 26540
rect 22796 26528 22802 26580
rect 23934 26528 23940 26580
rect 23992 26568 23998 26580
rect 25774 26568 25780 26580
rect 23992 26540 24992 26568
rect 25735 26540 25780 26568
rect 23992 26528 23998 26540
rect 15565 26503 15623 26509
rect 15565 26500 15577 26503
rect 12406 26472 15577 26500
rect 12406 26432 12434 26472
rect 15565 26469 15577 26472
rect 15611 26469 15623 26503
rect 19150 26500 19156 26512
rect 15565 26463 15623 26469
rect 15672 26472 19156 26500
rect 12618 26432 12624 26444
rect 11164 26404 12434 26432
rect 12531 26404 12624 26432
rect 10778 26364 10784 26376
rect 9640 26336 9996 26364
rect 10739 26336 10784 26364
rect 9640 26324 9646 26336
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 10870 26324 10876 26376
rect 10928 26364 10934 26376
rect 11974 26364 11980 26376
rect 10928 26336 10973 26364
rect 11935 26336 11980 26364
rect 10928 26324 10934 26336
rect 11974 26324 11980 26336
rect 12032 26324 12038 26376
rect 12158 26324 12164 26376
rect 12216 26364 12222 26376
rect 12544 26364 12572 26404
rect 12618 26392 12624 26404
rect 12676 26432 12682 26444
rect 14553 26435 14611 26441
rect 14553 26432 14565 26435
rect 12676 26404 14565 26432
rect 12676 26392 12682 26404
rect 14553 26401 14565 26404
rect 14599 26401 14611 26435
rect 14553 26395 14611 26401
rect 14274 26364 14280 26376
rect 12216 26336 12572 26364
rect 14235 26336 14280 26364
rect 12216 26324 12222 26336
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 15672 26364 15700 26472
rect 19150 26460 19156 26472
rect 19208 26460 19214 26512
rect 19705 26503 19763 26509
rect 19705 26469 19717 26503
rect 19751 26500 19763 26503
rect 20622 26500 20628 26512
rect 19751 26472 20628 26500
rect 19751 26469 19763 26472
rect 19705 26463 19763 26469
rect 20622 26460 20628 26472
rect 20680 26460 20686 26512
rect 24857 26503 24915 26509
rect 24857 26469 24869 26503
rect 24903 26469 24915 26503
rect 24857 26463 24915 26469
rect 15930 26432 15936 26444
rect 15891 26404 15936 26432
rect 15930 26392 15936 26404
rect 15988 26392 15994 26444
rect 16025 26435 16083 26441
rect 16025 26401 16037 26435
rect 16071 26432 16083 26435
rect 16114 26432 16120 26444
rect 16071 26404 16120 26432
rect 16071 26401 16083 26404
rect 16025 26395 16083 26401
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 24872 26432 24900 26463
rect 23492 26404 24900 26432
rect 24964 26432 24992 26540
rect 25774 26528 25780 26540
rect 25832 26528 25838 26580
rect 26145 26571 26203 26577
rect 26145 26537 26157 26571
rect 26191 26568 26203 26571
rect 26605 26571 26663 26577
rect 26605 26568 26617 26571
rect 26191 26540 26617 26568
rect 26191 26537 26203 26540
rect 26145 26531 26203 26537
rect 26605 26537 26617 26540
rect 26651 26537 26663 26571
rect 26786 26568 26792 26580
rect 26747 26540 26792 26568
rect 26605 26531 26663 26537
rect 26786 26528 26792 26540
rect 26844 26528 26850 26580
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 27798 26568 27804 26580
rect 27488 26540 27804 26568
rect 27488 26528 27494 26540
rect 27798 26528 27804 26540
rect 27856 26528 27862 26580
rect 27982 26568 27988 26580
rect 27943 26540 27988 26568
rect 27982 26528 27988 26540
rect 28040 26528 28046 26580
rect 30282 26568 30288 26580
rect 28092 26540 30288 26568
rect 27614 26460 27620 26512
rect 27672 26500 27678 26512
rect 28000 26500 28028 26528
rect 27672 26472 28028 26500
rect 27672 26460 27678 26472
rect 26053 26435 26111 26441
rect 26053 26432 26065 26435
rect 24964 26404 26065 26432
rect 15580 26336 15700 26364
rect 15749 26367 15807 26373
rect 8570 26296 8576 26308
rect 8312 26268 8576 26296
rect 8570 26256 8576 26268
rect 8628 26296 8634 26308
rect 9122 26296 9128 26308
rect 8628 26268 9128 26296
rect 8628 26256 8634 26268
rect 9122 26256 9128 26268
rect 9180 26256 9186 26308
rect 11054 26296 11060 26308
rect 11015 26268 11060 26296
rect 11054 26256 11060 26268
rect 11112 26256 11118 26308
rect 12069 26299 12127 26305
rect 12069 26265 12081 26299
rect 12115 26296 12127 26299
rect 12773 26299 12831 26305
rect 12773 26296 12785 26299
rect 12115 26268 12785 26296
rect 12115 26265 12127 26268
rect 12069 26259 12127 26265
rect 12773 26265 12785 26268
rect 12819 26265 12831 26299
rect 12773 26259 12831 26265
rect 12989 26299 13047 26305
rect 12989 26265 13001 26299
rect 13035 26296 13047 26299
rect 15580 26296 15608 26336
rect 15749 26333 15761 26367
rect 15795 26333 15807 26367
rect 15749 26327 15807 26333
rect 13035 26268 15608 26296
rect 13035 26265 13047 26268
rect 12989 26259 13047 26265
rect 15764 26240 15792 26327
rect 15838 26324 15844 26376
rect 15896 26364 15902 26376
rect 17586 26364 17592 26376
rect 15896 26336 17592 26364
rect 15896 26324 15902 26336
rect 17586 26324 17592 26336
rect 17644 26324 17650 26376
rect 17865 26367 17923 26373
rect 17865 26333 17877 26367
rect 17911 26364 17923 26367
rect 18598 26364 18604 26376
rect 17911 26336 18604 26364
rect 17911 26333 17923 26336
rect 17865 26327 17923 26333
rect 18598 26324 18604 26336
rect 18656 26324 18662 26376
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 20254 26364 20260 26376
rect 19475 26336 20260 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 20254 26324 20260 26336
rect 20312 26324 20318 26376
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21177 26367 21235 26373
rect 21177 26364 21189 26367
rect 20956 26336 21189 26364
rect 20956 26324 20962 26336
rect 21177 26333 21189 26336
rect 21223 26364 21235 26367
rect 21818 26364 21824 26376
rect 21223 26336 21824 26364
rect 21223 26333 21235 26336
rect 21177 26327 21235 26333
rect 21818 26324 21824 26336
rect 21876 26324 21882 26376
rect 19705 26299 19763 26305
rect 19705 26265 19717 26299
rect 19751 26296 19763 26299
rect 19978 26296 19984 26308
rect 19751 26268 19984 26296
rect 19751 26265 19763 26268
rect 19705 26259 19763 26265
rect 19978 26256 19984 26268
rect 20036 26256 20042 26308
rect 21444 26299 21502 26305
rect 21444 26265 21456 26299
rect 21490 26296 21502 26299
rect 23492 26296 23520 26404
rect 26053 26401 26065 26404
rect 26099 26401 26111 26435
rect 28092 26432 28120 26540
rect 30282 26528 30288 26540
rect 30340 26528 30346 26580
rect 29825 26503 29883 26509
rect 29825 26469 29837 26503
rect 29871 26500 29883 26503
rect 33870 26500 33876 26512
rect 29871 26472 33876 26500
rect 29871 26469 29883 26472
rect 29825 26463 29883 26469
rect 26053 26395 26111 26401
rect 27724 26404 28120 26432
rect 23566 26324 23572 26376
rect 23624 26364 23630 26376
rect 23753 26367 23811 26373
rect 23753 26364 23765 26367
rect 23624 26336 23765 26364
rect 23624 26324 23630 26336
rect 23753 26333 23765 26336
rect 23799 26333 23811 26367
rect 24026 26364 24032 26376
rect 23987 26336 24032 26364
rect 23753 26327 23811 26333
rect 24026 26324 24032 26336
rect 24084 26324 24090 26376
rect 24302 26324 24308 26376
rect 24360 26364 24366 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24360 26336 24593 26364
rect 24360 26324 24366 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24670 26324 24676 26376
rect 24728 26364 24734 26376
rect 24728 26336 24773 26364
rect 24728 26324 24734 26336
rect 26142 26324 26148 26376
rect 26200 26364 26206 26376
rect 26200 26336 26245 26364
rect 26200 26324 26206 26336
rect 27338 26324 27344 26376
rect 27396 26364 27402 26376
rect 27724 26373 27752 26404
rect 27709 26367 27767 26373
rect 27709 26364 27721 26367
rect 27396 26336 27721 26364
rect 27396 26324 27402 26336
rect 27709 26333 27721 26336
rect 27755 26333 27767 26367
rect 27890 26364 27896 26376
rect 27851 26336 27896 26364
rect 27709 26327 27767 26333
rect 27890 26324 27896 26336
rect 27948 26324 27954 26376
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26364 28227 26367
rect 28258 26364 28264 26376
rect 28215 26336 28264 26364
rect 28215 26333 28227 26336
rect 28169 26327 28227 26333
rect 28258 26324 28264 26336
rect 28316 26364 28322 26376
rect 28626 26364 28632 26376
rect 28316 26336 28632 26364
rect 28316 26324 28322 26336
rect 28626 26324 28632 26336
rect 28684 26324 28690 26376
rect 28994 26364 29000 26376
rect 28955 26336 29000 26364
rect 28994 26324 29000 26336
rect 29052 26324 29058 26376
rect 29181 26367 29239 26373
rect 29181 26333 29193 26367
rect 29227 26364 29239 26367
rect 29840 26364 29868 26463
rect 33870 26460 33876 26472
rect 33928 26460 33934 26512
rect 29227 26336 29868 26364
rect 30009 26367 30067 26373
rect 29227 26333 29239 26336
rect 29181 26327 29239 26333
rect 30009 26333 30021 26367
rect 30055 26364 30067 26367
rect 33594 26364 33600 26376
rect 30055 26336 33600 26364
rect 30055 26333 30067 26336
rect 30009 26327 30067 26333
rect 21490 26268 23520 26296
rect 24857 26299 24915 26305
rect 21490 26265 21502 26268
rect 21444 26259 21502 26265
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 24946 26296 24952 26308
rect 24903 26268 24952 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 24946 26256 24952 26268
rect 25004 26256 25010 26308
rect 26326 26256 26332 26308
rect 26384 26296 26390 26308
rect 26973 26299 27031 26305
rect 26973 26296 26985 26299
rect 26384 26268 26985 26296
rect 26384 26256 26390 26268
rect 26973 26265 26985 26268
rect 27019 26265 27031 26299
rect 26973 26259 27031 26265
rect 29730 26256 29736 26308
rect 29788 26296 29794 26308
rect 30024 26296 30052 26327
rect 33594 26324 33600 26336
rect 33652 26324 33658 26376
rect 29788 26268 30052 26296
rect 29788 26256 29794 26268
rect 12621 26231 12679 26237
rect 12621 26197 12633 26231
rect 12667 26228 12679 26231
rect 12894 26228 12900 26240
rect 12667 26200 12900 26228
rect 12667 26197 12679 26200
rect 12621 26191 12679 26197
rect 12894 26188 12900 26200
rect 12952 26188 12958 26240
rect 15746 26188 15752 26240
rect 15804 26188 15810 26240
rect 17402 26188 17408 26240
rect 17460 26228 17466 26240
rect 17773 26231 17831 26237
rect 17773 26228 17785 26231
rect 17460 26200 17785 26228
rect 17460 26188 17466 26200
rect 17773 26197 17785 26200
rect 17819 26228 17831 26231
rect 19426 26228 19432 26240
rect 17819 26200 19432 26228
rect 17819 26197 17831 26200
rect 17773 26191 17831 26197
rect 19426 26188 19432 26200
rect 19484 26228 19490 26240
rect 19521 26231 19579 26237
rect 19521 26228 19533 26231
rect 19484 26200 19533 26228
rect 19484 26188 19490 26200
rect 19521 26197 19533 26200
rect 19567 26197 19579 26231
rect 19521 26191 19579 26197
rect 26234 26188 26240 26240
rect 26292 26228 26298 26240
rect 26763 26231 26821 26237
rect 26763 26228 26775 26231
rect 26292 26200 26775 26228
rect 26292 26188 26298 26200
rect 26763 26197 26775 26200
rect 26809 26197 26821 26231
rect 26763 26191 26821 26197
rect 27062 26188 27068 26240
rect 27120 26228 27126 26240
rect 27433 26231 27491 26237
rect 27433 26228 27445 26231
rect 27120 26200 27445 26228
rect 27120 26188 27126 26200
rect 27433 26197 27445 26200
rect 27479 26197 27491 26231
rect 29086 26228 29092 26240
rect 29047 26200 29092 26228
rect 27433 26191 27491 26197
rect 29086 26188 29092 26200
rect 29144 26188 29150 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 8573 26027 8631 26033
rect 8573 25993 8585 26027
rect 8619 26024 8631 26027
rect 8846 26024 8852 26036
rect 8619 25996 8852 26024
rect 8619 25993 8631 25996
rect 8573 25987 8631 25993
rect 8846 25984 8852 25996
rect 8904 25984 8910 26036
rect 11054 25984 11060 26036
rect 11112 26024 11118 26036
rect 11793 26027 11851 26033
rect 11793 26024 11805 26027
rect 11112 25996 11805 26024
rect 11112 25984 11118 25996
rect 11793 25993 11805 25996
rect 11839 25993 11851 26027
rect 12710 26024 12716 26036
rect 11793 25987 11851 25993
rect 12360 25996 12716 26024
rect 8754 25956 8760 25968
rect 8715 25928 8760 25956
rect 8754 25916 8760 25928
rect 8812 25916 8818 25968
rect 8941 25959 8999 25965
rect 8941 25925 8953 25959
rect 8987 25956 8999 25959
rect 9493 25959 9551 25965
rect 9493 25956 9505 25959
rect 8987 25928 9505 25956
rect 8987 25925 8999 25928
rect 8941 25919 8999 25925
rect 9493 25925 9505 25928
rect 9539 25925 9551 25959
rect 12360 25956 12388 25996
rect 12710 25984 12716 25996
rect 12768 25984 12774 26036
rect 13817 26027 13875 26033
rect 13817 25993 13829 26027
rect 13863 26024 13875 26027
rect 14274 26024 14280 26036
rect 13863 25996 14280 26024
rect 13863 25993 13875 25996
rect 13817 25987 13875 25993
rect 14274 25984 14280 25996
rect 14332 25984 14338 26036
rect 15841 26027 15899 26033
rect 15841 25993 15853 26027
rect 15887 26024 15899 26027
rect 15930 26024 15936 26036
rect 15887 25996 15936 26024
rect 15887 25993 15899 25996
rect 15841 25987 15899 25993
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 17218 26024 17224 26036
rect 17179 25996 17224 26024
rect 17218 25984 17224 25996
rect 17276 25984 17282 26036
rect 17389 26027 17447 26033
rect 17389 25993 17401 26027
rect 17435 26024 17447 26027
rect 25685 26027 25743 26033
rect 17435 25996 18184 26024
rect 17435 25993 17447 25996
rect 17389 25987 17447 25993
rect 17586 25956 17592 25968
rect 9493 25919 9551 25925
rect 11716 25928 12388 25956
rect 17547 25928 17592 25956
rect 9306 25848 9312 25900
rect 9364 25888 9370 25900
rect 9401 25891 9459 25897
rect 9401 25888 9413 25891
rect 9364 25860 9413 25888
rect 9364 25848 9370 25860
rect 9401 25857 9413 25860
rect 9447 25857 9459 25891
rect 9582 25888 9588 25900
rect 9543 25860 9588 25888
rect 9401 25851 9459 25857
rect 9582 25848 9588 25860
rect 9640 25848 9646 25900
rect 11716 25897 11744 25928
rect 17586 25916 17592 25928
rect 17644 25916 17650 25968
rect 18046 25916 18052 25968
rect 18104 25956 18110 25968
rect 18156 25965 18184 25996
rect 25685 25993 25697 26027
rect 25731 26024 25743 26027
rect 26326 26024 26332 26036
rect 25731 25996 26332 26024
rect 25731 25993 25743 25996
rect 25685 25987 25743 25993
rect 26326 25984 26332 25996
rect 26384 25984 26390 26036
rect 27522 25984 27528 26036
rect 27580 26024 27586 26036
rect 27580 25996 27752 26024
rect 27580 25984 27586 25996
rect 18141 25959 18199 25965
rect 18141 25956 18153 25959
rect 18104 25928 18153 25956
rect 18104 25916 18110 25928
rect 18141 25925 18153 25928
rect 18187 25925 18199 25959
rect 18141 25919 18199 25925
rect 20622 25916 20628 25968
rect 20680 25965 20686 25968
rect 20680 25956 20692 25965
rect 25869 25959 25927 25965
rect 20680 25928 20725 25956
rect 20680 25919 20692 25928
rect 25869 25925 25881 25959
rect 25915 25956 25927 25959
rect 26234 25956 26240 25968
rect 25915 25928 26240 25956
rect 25915 25925 25927 25928
rect 25869 25919 25927 25925
rect 20680 25916 20686 25919
rect 26234 25916 26240 25928
rect 26292 25956 26298 25968
rect 27614 25956 27620 25968
rect 26292 25928 26464 25956
rect 26292 25916 26298 25928
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11790 25848 11796 25900
rect 11848 25888 11854 25900
rect 11885 25891 11943 25897
rect 11885 25888 11897 25891
rect 11848 25860 11897 25888
rect 11848 25848 11854 25860
rect 11885 25857 11897 25860
rect 11931 25857 11943 25891
rect 11885 25851 11943 25857
rect 12434 25848 12440 25900
rect 12492 25888 12498 25900
rect 12710 25897 12716 25900
rect 12492 25860 12537 25888
rect 12492 25848 12498 25860
rect 12704 25851 12716 25897
rect 12768 25888 12774 25900
rect 15749 25891 15807 25897
rect 12768 25860 12804 25888
rect 12710 25848 12716 25851
rect 12768 25848 12774 25860
rect 15749 25857 15761 25891
rect 15795 25888 15807 25891
rect 15838 25888 15844 25900
rect 15795 25860 15844 25888
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 15838 25848 15844 25860
rect 15896 25848 15902 25900
rect 20898 25888 20904 25900
rect 20859 25860 20904 25888
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 22646 25848 22652 25900
rect 22704 25888 22710 25900
rect 23382 25888 23388 25900
rect 22704 25860 23388 25888
rect 22704 25848 22710 25860
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 26436 25897 26464 25928
rect 27448 25928 27620 25956
rect 27448 25897 27476 25928
rect 27614 25916 27620 25928
rect 27672 25916 27678 25968
rect 27724 25897 27752 25996
rect 28988 25959 29046 25965
rect 28988 25925 29000 25959
rect 29034 25956 29046 25959
rect 29086 25956 29092 25968
rect 29034 25928 29092 25956
rect 29034 25925 29046 25928
rect 28988 25919 29046 25925
rect 29086 25916 29092 25928
rect 29144 25916 29150 25968
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 26421 25891 26479 25897
rect 26421 25857 26433 25891
rect 26467 25857 26479 25891
rect 26421 25851 26479 25857
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27525 25891 27583 25897
rect 27525 25857 27537 25891
rect 27571 25857 27583 25891
rect 27525 25851 27583 25857
rect 27709 25891 27767 25897
rect 27709 25857 27721 25891
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 14829 25823 14887 25829
rect 14829 25789 14841 25823
rect 14875 25820 14887 25823
rect 15194 25820 15200 25832
rect 14875 25792 15200 25820
rect 14875 25789 14887 25792
rect 14829 25783 14887 25789
rect 15194 25780 15200 25792
rect 15252 25780 15258 25832
rect 15289 25823 15347 25829
rect 15289 25789 15301 25823
rect 15335 25820 15347 25823
rect 16114 25820 16120 25832
rect 15335 25792 16120 25820
rect 15335 25789 15347 25792
rect 15289 25783 15347 25789
rect 16114 25780 16120 25792
rect 16172 25780 16178 25832
rect 25608 25820 25636 25851
rect 26326 25820 26332 25832
rect 25608 25792 26332 25820
rect 26326 25780 26332 25792
rect 26384 25820 26390 25832
rect 26786 25820 26792 25832
rect 26384 25792 26792 25820
rect 26384 25780 26390 25792
rect 26786 25780 26792 25792
rect 26844 25780 26850 25832
rect 27540 25820 27568 25851
rect 27798 25848 27804 25900
rect 27856 25888 27862 25900
rect 27856 25860 27901 25888
rect 27856 25848 27862 25860
rect 28258 25848 28264 25900
rect 28316 25888 28322 25900
rect 30742 25888 30748 25900
rect 28316 25860 30144 25888
rect 30703 25860 30748 25888
rect 28316 25848 28322 25860
rect 27614 25820 27620 25832
rect 27527 25792 27620 25820
rect 27614 25780 27620 25792
rect 27672 25820 27678 25832
rect 28074 25820 28080 25832
rect 27672 25792 28080 25820
rect 27672 25780 27678 25792
rect 28074 25780 28080 25792
rect 28132 25780 28138 25832
rect 28721 25823 28779 25829
rect 28721 25789 28733 25823
rect 28767 25789 28779 25823
rect 28721 25783 28779 25789
rect 30116 25820 30144 25860
rect 30742 25848 30748 25860
rect 30800 25848 30806 25900
rect 37461 25891 37519 25897
rect 37461 25857 37473 25891
rect 37507 25888 37519 25891
rect 38378 25888 38384 25900
rect 37507 25860 38384 25888
rect 37507 25857 37519 25860
rect 37461 25851 37519 25857
rect 38378 25848 38384 25860
rect 38436 25848 38442 25900
rect 30653 25823 30711 25829
rect 30653 25820 30665 25823
rect 30116 25792 30665 25820
rect 14274 25712 14280 25764
rect 14332 25752 14338 25764
rect 14918 25752 14924 25764
rect 14332 25724 14924 25752
rect 14332 25712 14338 25724
rect 14918 25712 14924 25724
rect 14976 25752 14982 25764
rect 15105 25755 15163 25761
rect 15105 25752 15117 25755
rect 14976 25724 15117 25752
rect 14976 25712 14982 25724
rect 15105 25721 15117 25724
rect 15151 25721 15163 25755
rect 15105 25715 15163 25721
rect 18325 25755 18383 25761
rect 18325 25721 18337 25755
rect 18371 25752 18383 25755
rect 18598 25752 18604 25764
rect 18371 25724 18604 25752
rect 18371 25721 18383 25724
rect 18325 25715 18383 25721
rect 18598 25712 18604 25724
rect 18656 25712 18662 25764
rect 21818 25712 21824 25764
rect 21876 25752 21882 25764
rect 24673 25755 24731 25761
rect 24673 25752 24685 25755
rect 21876 25724 24685 25752
rect 21876 25712 21882 25724
rect 24673 25721 24685 25724
rect 24719 25752 24731 25755
rect 25222 25752 25228 25764
rect 24719 25724 25228 25752
rect 24719 25721 24731 25724
rect 24673 25715 24731 25721
rect 25222 25712 25228 25724
rect 25280 25752 25286 25764
rect 28736 25752 28764 25783
rect 30116 25761 30144 25792
rect 30653 25789 30665 25792
rect 30699 25789 30711 25823
rect 30653 25783 30711 25789
rect 25280 25724 28764 25752
rect 30101 25755 30159 25761
rect 25280 25712 25286 25724
rect 30101 25721 30113 25755
rect 30147 25721 30159 25755
rect 30101 25715 30159 25721
rect 17402 25684 17408 25696
rect 17363 25656 17408 25684
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 19521 25687 19579 25693
rect 19521 25684 19533 25687
rect 19484 25656 19533 25684
rect 19484 25644 19490 25656
rect 19521 25653 19533 25656
rect 19567 25684 19579 25687
rect 19886 25684 19892 25696
rect 19567 25656 19892 25684
rect 19567 25653 19579 25656
rect 19521 25647 19579 25653
rect 19886 25644 19892 25656
rect 19944 25644 19950 25696
rect 25869 25687 25927 25693
rect 25869 25653 25881 25687
rect 25915 25684 25927 25687
rect 26142 25684 26148 25696
rect 25915 25656 26148 25684
rect 25915 25653 25927 25656
rect 25869 25647 25927 25653
rect 26142 25644 26148 25656
rect 26200 25644 26206 25696
rect 26510 25684 26516 25696
rect 26471 25656 26516 25684
rect 26510 25644 26516 25656
rect 26568 25644 26574 25696
rect 26602 25644 26608 25696
rect 26660 25684 26666 25696
rect 27249 25687 27307 25693
rect 27249 25684 27261 25687
rect 26660 25656 27261 25684
rect 26660 25644 26666 25656
rect 27249 25653 27261 25656
rect 27295 25653 27307 25687
rect 27249 25647 27307 25653
rect 31113 25687 31171 25693
rect 31113 25653 31125 25687
rect 31159 25684 31171 25687
rect 31386 25684 31392 25696
rect 31159 25656 31392 25684
rect 31159 25653 31171 25656
rect 31113 25647 31171 25653
rect 31386 25644 31392 25656
rect 31444 25644 31450 25696
rect 37553 25687 37611 25693
rect 37553 25653 37565 25687
rect 37599 25684 37611 25687
rect 38102 25684 38108 25696
rect 37599 25656 38108 25684
rect 37599 25653 37611 25656
rect 37553 25647 37611 25653
rect 38102 25644 38108 25656
rect 38160 25644 38166 25696
rect 38286 25684 38292 25696
rect 38247 25656 38292 25684
rect 38286 25644 38292 25656
rect 38344 25644 38350 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 4062 25480 4068 25492
rect 4023 25452 4068 25480
rect 4062 25440 4068 25452
rect 4120 25440 4126 25492
rect 12710 25480 12716 25492
rect 12671 25452 12716 25480
rect 12710 25440 12716 25452
rect 12768 25440 12774 25492
rect 14918 25480 14924 25492
rect 14879 25452 14924 25480
rect 14918 25440 14924 25452
rect 14976 25440 14982 25492
rect 15289 25483 15347 25489
rect 15289 25449 15301 25483
rect 15335 25480 15347 25483
rect 15746 25480 15752 25492
rect 15335 25452 15752 25480
rect 15335 25449 15347 25452
rect 15289 25443 15347 25449
rect 15746 25440 15752 25452
rect 15804 25440 15810 25492
rect 18046 25480 18052 25492
rect 18007 25452 18052 25480
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 19705 25483 19763 25489
rect 19705 25449 19717 25483
rect 19751 25480 19763 25483
rect 19978 25480 19984 25492
rect 19751 25452 19984 25480
rect 19751 25449 19763 25452
rect 19705 25443 19763 25449
rect 19978 25440 19984 25452
rect 20036 25440 20042 25492
rect 23753 25483 23811 25489
rect 23753 25449 23765 25483
rect 23799 25480 23811 25483
rect 24026 25480 24032 25492
rect 23799 25452 24032 25480
rect 23799 25449 23811 25452
rect 23753 25443 23811 25449
rect 24026 25440 24032 25452
rect 24084 25440 24090 25492
rect 24578 25480 24584 25492
rect 24539 25452 24584 25480
rect 24578 25440 24584 25452
rect 24636 25440 24642 25492
rect 27706 25480 27712 25492
rect 27448 25452 27712 25480
rect 24762 25372 24768 25424
rect 24820 25412 24826 25424
rect 27448 25412 27476 25452
rect 27706 25440 27712 25452
rect 27764 25480 27770 25492
rect 30374 25480 30380 25492
rect 27764 25452 30380 25480
rect 27764 25440 27770 25452
rect 30374 25440 30380 25452
rect 30432 25440 30438 25492
rect 24820 25384 27476 25412
rect 27525 25415 27583 25421
rect 24820 25372 24826 25384
rect 27525 25381 27537 25415
rect 27571 25412 27583 25415
rect 31846 25412 31852 25424
rect 27571 25384 31852 25412
rect 27571 25381 27583 25384
rect 27525 25375 27583 25381
rect 31846 25372 31852 25384
rect 31904 25372 31910 25424
rect 15930 25304 15936 25356
rect 15988 25344 15994 25356
rect 17126 25344 17132 25356
rect 15988 25316 17132 25344
rect 15988 25304 15994 25316
rect 17126 25304 17132 25316
rect 17184 25344 17190 25356
rect 18506 25344 18512 25356
rect 17184 25316 18512 25344
rect 17184 25304 17190 25316
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 19150 25304 19156 25356
rect 19208 25344 19214 25356
rect 19426 25344 19432 25356
rect 19208 25316 19432 25344
rect 19208 25304 19214 25316
rect 19426 25304 19432 25316
rect 19484 25344 19490 25356
rect 19613 25347 19671 25353
rect 19613 25344 19625 25347
rect 19484 25316 19625 25344
rect 19484 25304 19490 25316
rect 19613 25313 19625 25316
rect 19659 25313 19671 25347
rect 19613 25307 19671 25313
rect 21818 25304 21824 25356
rect 21876 25344 21882 25356
rect 22373 25347 22431 25353
rect 22373 25344 22385 25347
rect 21876 25316 22385 25344
rect 21876 25304 21882 25316
rect 22373 25313 22385 25316
rect 22419 25313 22431 25347
rect 22373 25307 22431 25313
rect 26510 25304 26516 25356
rect 26568 25344 26574 25356
rect 27341 25347 27399 25353
rect 27341 25344 27353 25347
rect 26568 25316 27353 25344
rect 26568 25304 26574 25316
rect 27341 25313 27353 25316
rect 27387 25313 27399 25347
rect 27341 25307 27399 25313
rect 30837 25347 30895 25353
rect 30837 25313 30849 25347
rect 30883 25344 30895 25347
rect 37826 25344 37832 25356
rect 30883 25316 31524 25344
rect 37787 25316 37832 25344
rect 30883 25313 30895 25316
rect 30837 25307 30895 25313
rect 31496 25288 31524 25316
rect 37826 25304 37832 25316
rect 37884 25304 37890 25356
rect 38102 25344 38108 25356
rect 38063 25316 38108 25344
rect 38102 25304 38108 25316
rect 38160 25304 38166 25356
rect 38286 25344 38292 25356
rect 38247 25316 38292 25344
rect 38286 25304 38292 25316
rect 38344 25304 38350 25356
rect 3878 25236 3884 25288
rect 3936 25276 3942 25288
rect 3973 25279 4031 25285
rect 3973 25276 3985 25279
rect 3936 25248 3985 25276
rect 3936 25236 3942 25248
rect 3973 25245 3985 25248
rect 4019 25245 4031 25279
rect 12894 25276 12900 25288
rect 12855 25248 12900 25276
rect 3973 25239 4031 25245
rect 12894 25236 12900 25248
rect 12952 25236 12958 25288
rect 14829 25279 14887 25285
rect 14829 25245 14841 25279
rect 14875 25276 14887 25279
rect 15194 25276 15200 25288
rect 14875 25248 15200 25276
rect 14875 25245 14887 25248
rect 14829 25239 14887 25245
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 17770 25236 17776 25288
rect 17828 25276 17834 25288
rect 18049 25279 18107 25285
rect 18049 25276 18061 25279
rect 17828 25248 18061 25276
rect 17828 25236 17834 25248
rect 18049 25245 18061 25248
rect 18095 25245 18107 25279
rect 18230 25276 18236 25288
rect 18191 25248 18236 25276
rect 18049 25239 18107 25245
rect 18230 25236 18236 25248
rect 18288 25236 18294 25288
rect 18598 25236 18604 25288
rect 18656 25276 18662 25288
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 18656 25248 19809 25276
rect 18656 25236 18662 25248
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 17126 25168 17132 25220
rect 17184 25208 17190 25220
rect 17221 25211 17279 25217
rect 17221 25208 17233 25211
rect 17184 25180 17233 25208
rect 17184 25168 17190 25180
rect 17221 25177 17233 25180
rect 17267 25177 17279 25211
rect 17221 25171 17279 25177
rect 17405 25211 17463 25217
rect 17405 25177 17417 25211
rect 17451 25208 17463 25211
rect 18414 25208 18420 25220
rect 17451 25180 18420 25208
rect 17451 25177 17463 25180
rect 17405 25171 17463 25177
rect 18414 25168 18420 25180
rect 18472 25168 18478 25220
rect 19812 25208 19840 25239
rect 19886 25236 19892 25288
rect 19944 25276 19950 25288
rect 19944 25248 19989 25276
rect 19944 25236 19950 25248
rect 20806 25236 20812 25288
rect 20864 25276 20870 25288
rect 21453 25279 21511 25285
rect 21453 25276 21465 25279
rect 20864 25248 21465 25276
rect 20864 25236 20870 25248
rect 21453 25245 21465 25248
rect 21499 25276 21511 25279
rect 22278 25276 22284 25288
rect 21499 25248 22284 25276
rect 21499 25245 21511 25248
rect 21453 25239 21511 25245
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 24762 25276 24768 25288
rect 24723 25248 24768 25276
rect 24762 25236 24768 25248
rect 24820 25236 24826 25288
rect 24857 25279 24915 25285
rect 24857 25245 24869 25279
rect 24903 25276 24915 25279
rect 26602 25276 26608 25288
rect 24903 25248 26608 25276
rect 24903 25245 24915 25248
rect 24857 25239 24915 25245
rect 26602 25236 26608 25248
rect 26660 25236 26666 25288
rect 27062 25276 27068 25288
rect 27023 25248 27068 25276
rect 27062 25236 27068 25248
rect 27120 25236 27126 25288
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 19812 25180 21404 25208
rect 16666 25100 16672 25152
rect 16724 25140 16730 25152
rect 17589 25143 17647 25149
rect 17589 25140 17601 25143
rect 16724 25112 17601 25140
rect 16724 25100 16730 25112
rect 17589 25109 17601 25112
rect 17635 25109 17647 25143
rect 21266 25140 21272 25152
rect 21227 25112 21272 25140
rect 17589 25103 17647 25109
rect 21266 25100 21272 25112
rect 21324 25100 21330 25152
rect 21376 25140 21404 25180
rect 22462 25168 22468 25220
rect 22520 25208 22526 25220
rect 22618 25211 22676 25217
rect 22618 25208 22630 25211
rect 22520 25180 22630 25208
rect 22520 25168 22526 25180
rect 22618 25177 22630 25180
rect 22664 25177 22676 25211
rect 22618 25171 22676 25177
rect 22830 25168 22836 25220
rect 22888 25208 22894 25220
rect 24581 25211 24639 25217
rect 24581 25208 24593 25211
rect 22888 25180 24593 25208
rect 22888 25168 22894 25180
rect 24581 25177 24593 25180
rect 24627 25177 24639 25211
rect 24581 25171 24639 25177
rect 26786 25168 26792 25220
rect 26844 25208 26850 25220
rect 27172 25208 27200 25239
rect 27246 25236 27252 25288
rect 27304 25276 27310 25288
rect 27304 25248 27844 25276
rect 27304 25236 27310 25248
rect 26844 25180 27200 25208
rect 27816 25208 27844 25248
rect 29086 25236 29092 25288
rect 29144 25276 29150 25288
rect 30561 25279 30619 25285
rect 30561 25276 30573 25279
rect 29144 25248 30573 25276
rect 29144 25236 29150 25248
rect 30561 25245 30573 25248
rect 30607 25245 30619 25279
rect 30561 25239 30619 25245
rect 30653 25279 30711 25285
rect 30653 25245 30665 25279
rect 30699 25276 30711 25279
rect 31297 25279 31355 25285
rect 31297 25276 31309 25279
rect 30699 25248 31309 25276
rect 30699 25245 30711 25248
rect 30653 25239 30711 25245
rect 31297 25245 31309 25248
rect 31343 25276 31355 25279
rect 31386 25276 31392 25288
rect 31343 25248 31392 25276
rect 31343 25245 31355 25248
rect 31297 25239 31355 25245
rect 31386 25236 31392 25248
rect 31444 25236 31450 25288
rect 31478 25236 31484 25288
rect 31536 25276 31542 25288
rect 31536 25248 31581 25276
rect 31536 25236 31542 25248
rect 27816 25180 30604 25208
rect 26844 25168 26850 25180
rect 23198 25140 23204 25152
rect 21376 25112 23204 25140
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 30576 25149 30604 25180
rect 30561 25143 30619 25149
rect 30561 25109 30573 25143
rect 30607 25109 30619 25143
rect 30561 25103 30619 25109
rect 30650 25100 30656 25152
rect 30708 25140 30714 25152
rect 31389 25143 31447 25149
rect 31389 25140 31401 25143
rect 30708 25112 31401 25140
rect 30708 25100 30714 25112
rect 31389 25109 31401 25112
rect 31435 25109 31447 25143
rect 31389 25103 31447 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 23198 24896 23204 24948
rect 23256 24936 23262 24948
rect 26326 24936 26332 24948
rect 23256 24908 25912 24936
rect 26287 24908 26332 24936
rect 23256 24896 23262 24908
rect 9398 24868 9404 24880
rect 9359 24840 9404 24868
rect 9398 24828 9404 24840
rect 9456 24828 9462 24880
rect 9766 24868 9772 24880
rect 9646 24843 9772 24868
rect 9631 24840 9772 24843
rect 9631 24837 9689 24840
rect 9631 24803 9643 24837
rect 9677 24803 9689 24837
rect 9766 24828 9772 24840
rect 9824 24828 9830 24880
rect 23658 24828 23664 24880
rect 23716 24868 23722 24880
rect 24673 24871 24731 24877
rect 24673 24868 24685 24871
rect 23716 24840 24685 24868
rect 23716 24828 23722 24840
rect 24673 24837 24685 24840
rect 24719 24837 24731 24871
rect 24673 24831 24731 24837
rect 24854 24828 24860 24880
rect 24912 24877 24918 24880
rect 25884 24877 25912 24908
rect 26326 24896 26332 24908
rect 26384 24896 26390 24948
rect 30009 24939 30067 24945
rect 30009 24905 30021 24939
rect 30055 24936 30067 24939
rect 30558 24936 30564 24948
rect 30055 24908 30564 24936
rect 30055 24905 30067 24908
rect 30009 24899 30067 24905
rect 30558 24896 30564 24908
rect 30616 24896 30622 24948
rect 31297 24939 31355 24945
rect 31297 24905 31309 24939
rect 31343 24936 31355 24939
rect 31478 24936 31484 24948
rect 31343 24908 31484 24936
rect 31343 24905 31355 24908
rect 31297 24899 31355 24905
rect 31478 24896 31484 24908
rect 31536 24896 31542 24948
rect 24912 24871 24931 24877
rect 24919 24837 24931 24871
rect 25869 24871 25927 24877
rect 24912 24831 24931 24837
rect 25639 24837 25697 24843
rect 24912 24828 24918 24831
rect 9631 24797 9689 24803
rect 10229 24803 10287 24809
rect 10229 24800 10241 24803
rect 9784 24772 10241 24800
rect 3881 24735 3939 24741
rect 3881 24701 3893 24735
rect 3927 24701 3939 24735
rect 4062 24732 4068 24744
rect 4023 24704 4068 24732
rect 3881 24695 3939 24701
rect 3896 24664 3924 24695
rect 4062 24692 4068 24704
rect 4120 24692 4126 24744
rect 5442 24732 5448 24744
rect 5403 24704 5448 24732
rect 5442 24692 5448 24704
rect 5500 24692 5506 24744
rect 4798 24664 4804 24676
rect 3896 24636 4804 24664
rect 4798 24624 4804 24636
rect 4856 24624 4862 24676
rect 9784 24673 9812 24772
rect 10229 24769 10241 24772
rect 10275 24769 10287 24803
rect 16022 24800 16028 24812
rect 15983 24772 16028 24800
rect 10229 24763 10287 24769
rect 16022 24760 16028 24772
rect 16080 24760 16086 24812
rect 17589 24803 17647 24809
rect 17589 24769 17601 24803
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24769 17831 24803
rect 17773 24763 17831 24769
rect 13722 24692 13728 24744
rect 13780 24732 13786 24744
rect 14185 24735 14243 24741
rect 14185 24732 14197 24735
rect 13780 24704 14197 24732
rect 13780 24692 13786 24704
rect 14185 24701 14197 24704
rect 14231 24701 14243 24735
rect 14366 24732 14372 24744
rect 14327 24704 14372 24732
rect 14185 24695 14243 24701
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 9769 24667 9827 24673
rect 9769 24633 9781 24667
rect 9815 24633 9827 24667
rect 17405 24667 17463 24673
rect 17405 24664 17417 24667
rect 9769 24627 9827 24633
rect 10244 24636 17417 24664
rect 8570 24556 8576 24608
rect 8628 24596 8634 24608
rect 9585 24599 9643 24605
rect 9585 24596 9597 24599
rect 8628 24568 9597 24596
rect 8628 24556 8634 24568
rect 9585 24565 9597 24568
rect 9631 24596 9643 24599
rect 10244 24596 10272 24636
rect 17405 24633 17417 24636
rect 17451 24633 17463 24667
rect 17405 24627 17463 24633
rect 10410 24596 10416 24608
rect 9631 24568 10272 24596
rect 10371 24568 10416 24596
rect 9631 24565 9643 24568
rect 9585 24559 9643 24565
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 17494 24556 17500 24608
rect 17552 24596 17558 24608
rect 17604 24596 17632 24763
rect 17788 24664 17816 24763
rect 17954 24760 17960 24812
rect 18012 24800 18018 24812
rect 18233 24803 18291 24809
rect 18233 24800 18245 24803
rect 18012 24772 18245 24800
rect 18012 24760 18018 24772
rect 18233 24769 18245 24772
rect 18279 24769 18291 24803
rect 18414 24800 18420 24812
rect 18375 24772 18420 24800
rect 18233 24763 18291 24769
rect 18414 24760 18420 24772
rect 18472 24800 18478 24812
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 18472 24772 19901 24800
rect 18472 24760 18478 24772
rect 19889 24769 19901 24772
rect 19935 24769 19947 24803
rect 20070 24800 20076 24812
rect 20031 24772 20076 24800
rect 19889 24763 19947 24769
rect 19904 24732 19932 24763
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20714 24800 20720 24812
rect 20675 24772 20720 24800
rect 20714 24760 20720 24772
rect 20772 24800 20778 24812
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 20772 24772 21189 24800
rect 20772 24760 20778 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 22830 24800 22836 24812
rect 21177 24763 21235 24769
rect 22066 24772 22836 24800
rect 20625 24735 20683 24741
rect 20625 24732 20637 24735
rect 19904 24704 20637 24732
rect 20625 24701 20637 24704
rect 20671 24732 20683 24735
rect 22066 24732 22094 24772
rect 22830 24760 22836 24772
rect 22888 24760 22894 24812
rect 25639 24803 25651 24837
rect 25685 24834 25697 24837
rect 25869 24837 25881 24871
rect 25915 24837 25927 24871
rect 26694 24868 26700 24880
rect 26607 24840 26700 24868
rect 25685 24806 25820 24834
rect 25869 24831 25927 24837
rect 25685 24803 25697 24806
rect 25639 24797 25697 24803
rect 25792 24800 25820 24806
rect 26510 24800 26516 24812
rect 25792 24772 26516 24800
rect 26510 24760 26516 24772
rect 26568 24760 26574 24812
rect 26620 24809 26648 24840
rect 26694 24828 26700 24840
rect 26752 24868 26758 24880
rect 27246 24868 27252 24880
rect 26752 24840 27252 24868
rect 26752 24828 26758 24840
rect 27246 24828 27252 24840
rect 27304 24828 27310 24880
rect 26605 24803 26663 24809
rect 26605 24769 26617 24803
rect 26651 24769 26663 24803
rect 27338 24800 27344 24812
rect 27299 24772 27344 24800
rect 26605 24763 26663 24769
rect 27338 24760 27344 24772
rect 27396 24760 27402 24812
rect 27525 24803 27583 24809
rect 27525 24769 27537 24803
rect 27571 24800 27583 24803
rect 27982 24800 27988 24812
rect 27571 24772 27988 24800
rect 27571 24769 27583 24772
rect 27525 24763 27583 24769
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 28074 24760 28080 24812
rect 28132 24800 28138 24812
rect 28261 24803 28319 24809
rect 28132 24772 28177 24800
rect 28132 24760 28138 24772
rect 28261 24769 28273 24803
rect 28307 24800 28319 24803
rect 28902 24800 28908 24812
rect 28307 24772 28908 24800
rect 28307 24769 28319 24772
rect 28261 24763 28319 24769
rect 28902 24760 28908 24772
rect 28960 24760 28966 24812
rect 29086 24800 29092 24812
rect 29047 24772 29092 24800
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 29273 24803 29331 24809
rect 29273 24769 29285 24803
rect 29319 24800 29331 24803
rect 29730 24800 29736 24812
rect 29319 24772 29736 24800
rect 29319 24769 29331 24772
rect 29273 24763 29331 24769
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 29950 24803 30008 24809
rect 29950 24800 29962 24803
rect 29840 24772 29962 24800
rect 20671 24704 22094 24732
rect 20671 24701 20683 24704
rect 20625 24695 20683 24701
rect 22278 24692 22284 24744
rect 22336 24732 22342 24744
rect 22557 24735 22615 24741
rect 22557 24732 22569 24735
rect 22336 24704 22569 24732
rect 22336 24692 22342 24704
rect 22557 24701 22569 24704
rect 22603 24701 22615 24735
rect 22557 24695 22615 24701
rect 26329 24735 26387 24741
rect 26329 24701 26341 24735
rect 26375 24732 26387 24735
rect 26786 24732 26792 24744
rect 26375 24704 26792 24732
rect 26375 24701 26387 24704
rect 26329 24695 26387 24701
rect 26786 24692 26792 24704
rect 26844 24692 26850 24744
rect 27614 24732 27620 24744
rect 27575 24704 27620 24732
rect 27614 24692 27620 24704
rect 27672 24692 27678 24744
rect 28166 24732 28172 24744
rect 28127 24704 28172 24732
rect 28166 24692 28172 24704
rect 28224 24692 28230 24744
rect 29840 24732 29868 24772
rect 29950 24769 29962 24772
rect 29996 24769 30008 24803
rect 29950 24763 30008 24769
rect 30469 24803 30527 24809
rect 30469 24769 30481 24803
rect 30515 24800 30527 24803
rect 30650 24800 30656 24812
rect 30515 24772 30656 24800
rect 30515 24769 30527 24772
rect 30469 24763 30527 24769
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 31110 24800 31116 24812
rect 31071 24772 31116 24800
rect 31110 24760 31116 24772
rect 31168 24760 31174 24812
rect 31386 24760 31392 24812
rect 31444 24800 31450 24812
rect 31444 24772 31489 24800
rect 31444 24760 31450 24772
rect 37274 24760 37280 24812
rect 37332 24800 37338 24812
rect 37461 24803 37519 24809
rect 37461 24800 37473 24803
rect 37332 24772 37473 24800
rect 37332 24760 37338 24772
rect 37461 24769 37473 24772
rect 37507 24769 37519 24803
rect 37461 24763 37519 24769
rect 30190 24732 30196 24744
rect 28920 24704 30196 24732
rect 20073 24667 20131 24673
rect 20073 24664 20085 24667
rect 17788 24636 20085 24664
rect 20073 24633 20085 24636
rect 20119 24664 20131 24667
rect 20346 24664 20352 24676
rect 20119 24636 20352 24664
rect 20119 24633 20131 24636
rect 20073 24627 20131 24633
rect 20346 24624 20352 24636
rect 20404 24624 20410 24676
rect 27632 24664 27660 24692
rect 28920 24664 28948 24704
rect 30190 24692 30196 24704
rect 30248 24692 30254 24744
rect 27632 24636 28948 24664
rect 28994 24624 29000 24676
rect 29052 24664 29058 24676
rect 29825 24667 29883 24673
rect 29825 24664 29837 24667
rect 29052 24636 29837 24664
rect 29052 24624 29058 24636
rect 29825 24633 29837 24636
rect 29871 24633 29883 24667
rect 29825 24627 29883 24633
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 17552 24568 18245 24596
rect 17552 24556 17558 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 21358 24596 21364 24608
rect 21319 24568 21364 24596
rect 18233 24559 18291 24565
rect 21358 24556 21364 24568
rect 21416 24556 21422 24608
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 24857 24599 24915 24605
rect 24857 24596 24869 24599
rect 24820 24568 24869 24596
rect 24820 24556 24826 24568
rect 24857 24565 24869 24568
rect 24903 24565 24915 24599
rect 24857 24559 24915 24565
rect 25041 24599 25099 24605
rect 25041 24565 25053 24599
rect 25087 24596 25099 24599
rect 25130 24596 25136 24608
rect 25087 24568 25136 24596
rect 25087 24565 25099 24568
rect 25041 24559 25099 24565
rect 25130 24556 25136 24568
rect 25188 24556 25194 24608
rect 25498 24596 25504 24608
rect 25459 24568 25504 24596
rect 25498 24556 25504 24568
rect 25556 24556 25562 24608
rect 25685 24599 25743 24605
rect 25685 24565 25697 24599
rect 25731 24596 25743 24599
rect 26326 24596 26332 24608
rect 25731 24568 26332 24596
rect 25731 24565 25743 24568
rect 25685 24559 25743 24565
rect 26326 24556 26332 24568
rect 26384 24556 26390 24608
rect 26513 24599 26571 24605
rect 26513 24565 26525 24599
rect 26559 24596 26571 24599
rect 26878 24596 26884 24608
rect 26559 24568 26884 24596
rect 26559 24565 26571 24568
rect 26513 24559 26571 24565
rect 26878 24556 26884 24568
rect 26936 24596 26942 24608
rect 27157 24599 27215 24605
rect 27157 24596 27169 24599
rect 26936 24568 27169 24596
rect 26936 24556 26942 24568
rect 27157 24565 27169 24568
rect 27203 24565 27215 24599
rect 27157 24559 27215 24565
rect 28626 24556 28632 24608
rect 28684 24596 28690 24608
rect 29181 24599 29239 24605
rect 29181 24596 29193 24599
rect 28684 24568 29193 24596
rect 28684 24556 28690 24568
rect 29181 24565 29193 24568
rect 29227 24565 29239 24599
rect 29181 24559 29239 24565
rect 30377 24599 30435 24605
rect 30377 24565 30389 24599
rect 30423 24596 30435 24599
rect 30929 24599 30987 24605
rect 30929 24596 30941 24599
rect 30423 24568 30941 24596
rect 30423 24565 30435 24568
rect 30377 24559 30435 24565
rect 30929 24565 30941 24568
rect 30975 24565 30987 24599
rect 30929 24559 30987 24565
rect 37553 24599 37611 24605
rect 37553 24565 37565 24599
rect 37599 24596 37611 24599
rect 38102 24596 38108 24608
rect 37599 24568 38108 24596
rect 37599 24565 37611 24568
rect 37553 24559 37611 24565
rect 38102 24556 38108 24568
rect 38160 24556 38166 24608
rect 38286 24596 38292 24608
rect 38247 24568 38292 24596
rect 38286 24556 38292 24568
rect 38344 24556 38350 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 4062 24392 4068 24404
rect 4023 24364 4068 24392
rect 4062 24352 4068 24364
rect 4120 24352 4126 24404
rect 9217 24395 9275 24401
rect 9217 24361 9229 24395
rect 9263 24392 9275 24395
rect 9398 24392 9404 24404
rect 9263 24364 9404 24392
rect 9263 24361 9275 24364
rect 9217 24355 9275 24361
rect 9398 24352 9404 24364
rect 9456 24352 9462 24404
rect 11701 24395 11759 24401
rect 11701 24361 11713 24395
rect 11747 24392 11759 24395
rect 11790 24392 11796 24404
rect 11747 24364 11796 24392
rect 11747 24361 11759 24364
rect 11701 24355 11759 24361
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 13722 24392 13728 24404
rect 13683 24364 13728 24392
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 14274 24352 14280 24404
rect 14332 24392 14338 24404
rect 19334 24392 19340 24404
rect 14332 24364 19340 24392
rect 14332 24352 14338 24364
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 22462 24392 22468 24404
rect 22423 24364 22468 24392
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 25041 24395 25099 24401
rect 25041 24361 25053 24395
rect 25087 24392 25099 24395
rect 25498 24392 25504 24404
rect 25087 24364 25504 24392
rect 25087 24361 25099 24364
rect 25041 24355 25099 24361
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 26510 24392 26516 24404
rect 26471 24364 26516 24392
rect 26510 24352 26516 24364
rect 26568 24352 26574 24404
rect 26694 24392 26700 24404
rect 26655 24364 26700 24392
rect 26694 24352 26700 24364
rect 26752 24352 26758 24404
rect 28902 24392 28908 24404
rect 28863 24364 28908 24392
rect 28902 24352 28908 24364
rect 28960 24352 28966 24404
rect 29730 24392 29736 24404
rect 29691 24364 29736 24392
rect 29730 24352 29736 24364
rect 29788 24352 29794 24404
rect 23661 24327 23719 24333
rect 23661 24324 23673 24327
rect 22946 24296 23673 24324
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 18693 24259 18751 24265
rect 18693 24256 18705 24259
rect 12584 24228 14872 24256
rect 12584 24216 12590 24228
rect 3878 24148 3884 24200
rect 3936 24188 3942 24200
rect 3973 24191 4031 24197
rect 3973 24188 3985 24191
rect 3936 24160 3985 24188
rect 3936 24148 3942 24160
rect 3973 24157 3985 24160
rect 4019 24157 4031 24191
rect 8570 24188 8576 24200
rect 8531 24160 8576 24188
rect 3973 24151 4031 24157
rect 8570 24148 8576 24160
rect 8628 24148 8634 24200
rect 9401 24191 9459 24197
rect 9401 24157 9413 24191
rect 9447 24188 9459 24191
rect 10226 24188 10232 24200
rect 9447 24160 10232 24188
rect 9447 24157 9459 24160
rect 9401 24151 9459 24157
rect 10226 24148 10232 24160
rect 10284 24148 10290 24200
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24188 10379 24191
rect 10367 24160 10732 24188
rect 10367 24157 10379 24160
rect 10321 24151 10379 24157
rect 10704 24132 10732 24160
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12989 24191 13047 24197
rect 12989 24188 13001 24191
rect 12400 24160 13001 24188
rect 12400 24148 12406 24160
rect 12989 24157 13001 24160
rect 13035 24157 13047 24191
rect 12989 24151 13047 24157
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 14090 24188 14096 24200
rect 13587 24160 14096 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24157 14795 24191
rect 14844 24188 14872 24228
rect 17328 24228 18705 24256
rect 16954 24191 17012 24197
rect 14844 24160 16804 24188
rect 14737 24151 14795 24157
rect 9585 24123 9643 24129
rect 9585 24089 9597 24123
rect 9631 24120 9643 24123
rect 10042 24120 10048 24132
rect 9631 24092 10048 24120
rect 9631 24089 9643 24092
rect 9585 24083 9643 24089
rect 10042 24080 10048 24092
rect 10100 24080 10106 24132
rect 10410 24080 10416 24132
rect 10468 24120 10474 24132
rect 10566 24123 10624 24129
rect 10566 24120 10578 24123
rect 10468 24092 10578 24120
rect 10468 24080 10474 24092
rect 10566 24089 10578 24092
rect 10612 24089 10624 24123
rect 10566 24083 10624 24089
rect 10686 24080 10692 24132
rect 10744 24120 10750 24132
rect 14752 24120 14780 24151
rect 10744 24092 14780 24120
rect 15004 24123 15062 24129
rect 10744 24080 10750 24092
rect 15004 24089 15016 24123
rect 15050 24120 15062 24123
rect 16666 24120 16672 24132
rect 15050 24092 16252 24120
rect 16627 24092 16672 24120
rect 15050 24089 15062 24092
rect 15004 24083 15062 24089
rect 8481 24055 8539 24061
rect 8481 24021 8493 24055
rect 8527 24052 8539 24055
rect 9030 24052 9036 24064
rect 8527 24024 9036 24052
rect 8527 24021 8539 24024
rect 8481 24015 8539 24021
rect 9030 24012 9036 24024
rect 9088 24012 9094 24064
rect 9122 24012 9128 24064
rect 9180 24052 9186 24064
rect 12897 24055 12955 24061
rect 12897 24052 12909 24055
rect 9180 24024 12909 24052
rect 9180 24012 9186 24024
rect 12897 24021 12909 24024
rect 12943 24052 12955 24055
rect 13354 24052 13360 24064
rect 12943 24024 13360 24052
rect 12943 24021 12955 24024
rect 12897 24015 12955 24021
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 15194 24012 15200 24064
rect 15252 24052 15258 24064
rect 16114 24052 16120 24064
rect 15252 24024 16120 24052
rect 15252 24012 15258 24024
rect 16114 24012 16120 24024
rect 16172 24012 16178 24064
rect 16224 24052 16252 24092
rect 16666 24080 16672 24092
rect 16724 24080 16730 24132
rect 16776 24120 16804 24160
rect 16954 24157 16966 24191
rect 17000 24188 17012 24191
rect 17328 24188 17356 24228
rect 17494 24188 17500 24200
rect 17000 24160 17356 24188
rect 17455 24160 17500 24188
rect 17000 24157 17012 24160
rect 16954 24151 17012 24157
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17696 24197 17724 24228
rect 18693 24225 18705 24228
rect 18739 24225 18751 24259
rect 22646 24256 22652 24268
rect 18693 24219 18751 24225
rect 21560 24228 22652 24256
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 17911 24191 17969 24197
rect 17911 24157 17923 24191
rect 17957 24188 17969 24191
rect 18506 24188 18512 24200
rect 17957 24160 18512 24188
rect 17957 24157 17969 24160
rect 17911 24151 17969 24157
rect 16776 24092 17080 24120
rect 16767 24055 16825 24061
rect 16767 24052 16779 24055
rect 16224 24024 16779 24052
rect 16767 24021 16779 24024
rect 16813 24021 16825 24055
rect 16767 24015 16825 24021
rect 16853 24055 16911 24061
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 16942 24052 16948 24064
rect 16899 24024 16948 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 17052 24052 17080 24092
rect 17586 24080 17592 24132
rect 17644 24120 17650 24132
rect 17788 24120 17816 24151
rect 18506 24148 18512 24160
rect 18564 24188 18570 24200
rect 18601 24191 18659 24197
rect 18601 24188 18613 24191
rect 18564 24160 18613 24188
rect 18564 24148 18570 24160
rect 18601 24157 18613 24160
rect 18647 24157 18659 24191
rect 18782 24188 18788 24200
rect 18743 24160 18788 24188
rect 18601 24151 18659 24157
rect 18782 24148 18788 24160
rect 18840 24188 18846 24200
rect 20070 24188 20076 24200
rect 18840 24160 20076 24188
rect 18840 24148 18846 24160
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20257 24123 20315 24129
rect 20257 24120 20269 24123
rect 17644 24092 17816 24120
rect 17972 24092 20269 24120
rect 17644 24080 17650 24092
rect 17972 24052 18000 24092
rect 20257 24089 20269 24092
rect 20303 24089 20315 24123
rect 20257 24083 20315 24089
rect 18138 24052 18144 24064
rect 17052 24024 18000 24052
rect 18099 24024 18144 24052
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 20806 24012 20812 24064
rect 20864 24052 20870 24064
rect 21560 24061 21588 24228
rect 22646 24216 22652 24228
rect 22704 24216 22710 24268
rect 22946 24197 22974 24296
rect 23661 24293 23673 24296
rect 23707 24293 23719 24327
rect 28074 24324 28080 24336
rect 23661 24287 23719 24293
rect 24872 24296 28080 24324
rect 24872 24256 24900 24296
rect 28074 24284 28080 24296
rect 28132 24284 28138 24336
rect 25130 24256 25136 24268
rect 23492 24228 24900 24256
rect 25091 24228 25136 24256
rect 22741 24191 22799 24197
rect 22741 24157 22753 24191
rect 22787 24157 22799 24191
rect 22741 24151 22799 24157
rect 22830 24188 22888 24194
rect 22830 24154 22842 24188
rect 22876 24154 22888 24188
rect 21545 24055 21603 24061
rect 21545 24052 21557 24055
rect 20864 24024 21557 24052
rect 20864 24012 20870 24024
rect 21545 24021 21557 24024
rect 21591 24021 21603 24055
rect 22756 24052 22784 24151
rect 22830 24148 22888 24154
rect 22930 24191 22988 24197
rect 22930 24157 22942 24191
rect 22976 24157 22988 24191
rect 22930 24151 22988 24157
rect 23106 24148 23112 24200
rect 23164 24188 23170 24200
rect 23492 24188 23520 24228
rect 23164 24160 23520 24188
rect 23569 24191 23627 24197
rect 23164 24148 23170 24160
rect 23569 24157 23581 24191
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 22845 24120 22873 24148
rect 23198 24120 23204 24132
rect 22845 24092 23204 24120
rect 23198 24080 23204 24092
rect 23256 24080 23262 24132
rect 23584 24064 23612 24151
rect 23750 24148 23756 24200
rect 23808 24188 23814 24200
rect 24872 24197 24900 24228
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 26786 24256 26792 24268
rect 26747 24228 26792 24256
rect 26786 24216 26792 24228
rect 26844 24216 26850 24268
rect 27801 24259 27859 24265
rect 27801 24225 27813 24259
rect 27847 24256 27859 24259
rect 28445 24259 28503 24265
rect 28445 24256 28457 24259
rect 27847 24228 28457 24256
rect 27847 24225 27859 24228
rect 27801 24219 27859 24225
rect 28445 24225 28457 24228
rect 28491 24225 28503 24259
rect 28626 24256 28632 24268
rect 28587 24228 28632 24256
rect 28445 24219 28503 24225
rect 28626 24216 28632 24228
rect 28684 24216 28690 24268
rect 30650 24256 30656 24268
rect 29932 24228 30656 24256
rect 24857 24191 24915 24197
rect 23808 24160 24808 24188
rect 23808 24148 23814 24160
rect 24780 24120 24808 24160
rect 24857 24157 24869 24191
rect 24903 24157 24915 24191
rect 24857 24151 24915 24157
rect 26878 24148 26884 24200
rect 26936 24188 26942 24200
rect 26936 24160 26981 24188
rect 26936 24148 26942 24160
rect 27338 24148 27344 24200
rect 27396 24188 27402 24200
rect 27709 24191 27767 24197
rect 27709 24188 27721 24191
rect 27396 24160 27721 24188
rect 27396 24148 27402 24160
rect 27709 24157 27721 24160
rect 27755 24157 27767 24191
rect 27709 24151 27767 24157
rect 27893 24191 27951 24197
rect 27893 24157 27905 24191
rect 27939 24188 27951 24191
rect 27982 24188 27988 24200
rect 27939 24160 27988 24188
rect 27939 24157 27951 24160
rect 27893 24151 27951 24157
rect 27982 24148 27988 24160
rect 28040 24148 28046 24200
rect 28258 24148 28264 24200
rect 28316 24188 28322 24200
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 28316 24160 28549 24188
rect 28316 24148 28322 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24188 28779 24191
rect 29178 24188 29184 24200
rect 28767 24160 29184 24188
rect 28767 24157 28779 24160
rect 28721 24151 28779 24157
rect 29178 24148 29184 24160
rect 29236 24148 29242 24200
rect 29932 24197 29960 24228
rect 30650 24216 30656 24228
rect 30708 24216 30714 24268
rect 37826 24256 37832 24268
rect 37787 24228 37832 24256
rect 37826 24216 37832 24228
rect 37884 24216 37890 24268
rect 38102 24256 38108 24268
rect 38063 24228 38108 24256
rect 38102 24216 38108 24228
rect 38160 24216 38166 24268
rect 38286 24256 38292 24268
rect 38247 24228 38292 24256
rect 38286 24216 38292 24228
rect 38344 24216 38350 24268
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 30190 24188 30196 24200
rect 30151 24160 30196 24188
rect 29917 24151 29975 24157
rect 30190 24148 30196 24160
rect 30248 24148 30254 24200
rect 27356 24120 27384 24148
rect 31110 24120 31116 24132
rect 24780 24092 27384 24120
rect 27448 24092 31116 24120
rect 23566 24052 23572 24064
rect 22756 24024 23572 24052
rect 21545 24015 21603 24021
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 24673 24055 24731 24061
rect 24673 24021 24685 24055
rect 24719 24052 24731 24055
rect 24762 24052 24768 24064
rect 24719 24024 24768 24052
rect 24719 24021 24731 24024
rect 24673 24015 24731 24021
rect 24762 24012 24768 24024
rect 24820 24012 24826 24064
rect 24854 24012 24860 24064
rect 24912 24052 24918 24064
rect 27448 24052 27476 24092
rect 31110 24080 31116 24092
rect 31168 24080 31174 24132
rect 24912 24024 27476 24052
rect 30101 24055 30159 24061
rect 24912 24012 24918 24024
rect 30101 24021 30113 24055
rect 30147 24052 30159 24055
rect 30282 24052 30288 24064
rect 30147 24024 30288 24052
rect 30147 24021 30159 24024
rect 30101 24015 30159 24021
rect 30282 24012 30288 24024
rect 30340 24012 30346 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 3878 23808 3884 23860
rect 3936 23848 3942 23860
rect 13814 23848 13820 23860
rect 3936 23820 13820 23848
rect 3936 23808 3942 23820
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 14090 23848 14096 23860
rect 14051 23820 14096 23848
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 16942 23848 16948 23860
rect 15396 23820 16948 23848
rect 10042 23789 10048 23792
rect 10029 23783 10048 23789
rect 10029 23749 10041 23783
rect 10029 23743 10048 23749
rect 10042 23740 10048 23743
rect 10100 23740 10106 23792
rect 10229 23783 10287 23789
rect 10229 23749 10241 23783
rect 10275 23749 10287 23783
rect 10229 23743 10287 23749
rect 9030 23712 9036 23724
rect 8991 23684 9036 23712
rect 9030 23672 9036 23684
rect 9088 23672 9094 23724
rect 9122 23672 9128 23724
rect 9180 23712 9186 23724
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 9180 23684 9229 23712
rect 9180 23672 9186 23684
rect 9217 23681 9229 23684
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23712 9459 23715
rect 9766 23712 9772 23724
rect 9447 23684 9772 23712
rect 9447 23681 9459 23684
rect 9401 23675 9459 23681
rect 9766 23672 9772 23684
rect 9824 23712 9830 23724
rect 10134 23712 10140 23724
rect 9824 23684 10140 23712
rect 9824 23672 9830 23684
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10244 23712 10272 23743
rect 11790 23740 11796 23792
rect 11848 23780 11854 23792
rect 12250 23780 12256 23792
rect 11848 23752 12256 23780
rect 11848 23740 11854 23752
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 15396 23780 15424 23820
rect 16942 23808 16948 23820
rect 17000 23808 17006 23860
rect 17586 23808 17592 23860
rect 17644 23848 17650 23860
rect 18782 23848 18788 23860
rect 17644 23820 18788 23848
rect 17644 23808 17650 23820
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 20441 23851 20499 23857
rect 20441 23817 20453 23851
rect 20487 23848 20499 23851
rect 20714 23848 20720 23860
rect 20487 23820 20720 23848
rect 20487 23817 20499 23820
rect 20441 23811 20499 23817
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 23934 23848 23940 23860
rect 22235 23820 23940 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 23934 23808 23940 23820
rect 23992 23808 23998 23860
rect 29178 23848 29184 23860
rect 29139 23820 29184 23848
rect 29178 23808 29184 23820
rect 29236 23808 29242 23860
rect 13280 23752 15424 23780
rect 12342 23712 12348 23724
rect 10244 23684 12348 23712
rect 12342 23672 12348 23684
rect 12400 23672 12406 23724
rect 13280 23721 13308 23752
rect 15470 23740 15476 23792
rect 15528 23780 15534 23792
rect 17313 23783 17371 23789
rect 17313 23780 17325 23783
rect 15528 23752 17325 23780
rect 15528 23740 15534 23752
rect 17313 23749 17325 23752
rect 17359 23749 17371 23783
rect 17313 23743 17371 23749
rect 18138 23740 18144 23792
rect 18196 23780 18202 23792
rect 19438 23783 19496 23789
rect 19438 23780 19450 23783
rect 18196 23752 19450 23780
rect 18196 23740 18202 23752
rect 19438 23749 19450 23752
rect 19484 23749 19496 23783
rect 20898 23780 20904 23792
rect 20859 23752 20904 23780
rect 19438 23743 19496 23749
rect 20898 23740 20904 23752
rect 20956 23740 20962 23792
rect 22278 23740 22284 23792
rect 22336 23780 22342 23792
rect 23569 23783 23627 23789
rect 23569 23780 23581 23783
rect 22336 23752 23581 23780
rect 22336 23740 22342 23752
rect 23569 23749 23581 23752
rect 23615 23749 23627 23783
rect 23569 23743 23627 23749
rect 23753 23783 23811 23789
rect 23753 23749 23765 23783
rect 23799 23780 23811 23783
rect 24946 23780 24952 23792
rect 23799 23752 24952 23780
rect 23799 23749 23811 23752
rect 23753 23743 23811 23749
rect 24946 23740 24952 23752
rect 25004 23780 25010 23792
rect 27798 23780 27804 23792
rect 25004 23752 27804 23780
rect 25004 23740 25010 23752
rect 27798 23740 27804 23752
rect 27856 23740 27862 23792
rect 29086 23740 29092 23792
rect 29144 23780 29150 23792
rect 29365 23783 29423 23789
rect 29365 23780 29377 23783
rect 29144 23752 29377 23780
rect 29144 23740 29150 23752
rect 29365 23749 29377 23752
rect 29411 23749 29423 23783
rect 29365 23743 29423 23749
rect 29549 23783 29607 23789
rect 29549 23749 29561 23783
rect 29595 23780 29607 23783
rect 29730 23780 29736 23792
rect 29595 23752 29736 23780
rect 29595 23749 29607 23752
rect 29549 23743 29607 23749
rect 29730 23740 29736 23752
rect 29788 23740 29794 23792
rect 35710 23780 35716 23792
rect 35671 23752 35716 23780
rect 35710 23740 35716 23752
rect 35768 23740 35774 23792
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23681 13323 23715
rect 13265 23675 13323 23681
rect 13354 23672 13360 23724
rect 13412 23712 13418 23724
rect 14274 23712 14280 23724
rect 13412 23684 13457 23712
rect 14235 23684 14280 23712
rect 13412 23672 13418 23684
rect 14274 23672 14280 23684
rect 14332 23672 14338 23724
rect 14737 23715 14795 23721
rect 14737 23681 14749 23715
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 13906 23644 13912 23656
rect 12483 23616 13912 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 13906 23604 13912 23616
rect 13964 23604 13970 23656
rect 14182 23604 14188 23656
rect 14240 23644 14246 23656
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 14240 23616 14381 23644
rect 14240 23604 14246 23616
rect 14369 23613 14381 23616
rect 14415 23613 14427 23647
rect 14752 23644 14780 23675
rect 15654 23672 15660 23724
rect 15712 23712 15718 23724
rect 17221 23715 17279 23721
rect 17221 23712 17233 23715
rect 15712 23684 17233 23712
rect 15712 23672 15718 23684
rect 17221 23681 17233 23684
rect 17267 23681 17279 23715
rect 17221 23675 17279 23681
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23712 17555 23715
rect 18414 23712 18420 23724
rect 17543 23684 18420 23712
rect 17543 23681 17555 23684
rect 17497 23675 17555 23681
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 22094 23672 22100 23724
rect 22152 23712 22158 23724
rect 24762 23721 24768 23724
rect 22833 23715 22891 23721
rect 22833 23712 22845 23715
rect 22152 23684 22845 23712
rect 22152 23672 22158 23684
rect 22833 23681 22845 23684
rect 22879 23681 22891 23715
rect 24756 23712 24768 23721
rect 24723 23684 24768 23712
rect 22833 23675 22891 23681
rect 24756 23675 24768 23684
rect 24762 23672 24768 23675
rect 24820 23672 24826 23724
rect 26970 23672 26976 23724
rect 27028 23712 27034 23724
rect 28353 23715 28411 23721
rect 28353 23712 28365 23715
rect 27028 23684 28365 23712
rect 27028 23672 27034 23684
rect 28353 23681 28365 23684
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 18138 23644 18144 23656
rect 14752 23616 18144 23644
rect 14369 23607 14427 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23644 19763 23647
rect 22186 23644 22192 23656
rect 19751 23616 20852 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 9033 23579 9091 23585
rect 9033 23545 9045 23579
rect 9079 23576 9091 23579
rect 10870 23576 10876 23588
rect 9079 23548 10876 23576
rect 9079 23545 9091 23548
rect 9033 23539 9091 23545
rect 10870 23536 10876 23548
rect 10928 23536 10934 23588
rect 13633 23579 13691 23585
rect 13633 23545 13645 23579
rect 13679 23576 13691 23579
rect 17497 23579 17555 23585
rect 13679 23548 14320 23576
rect 13679 23545 13691 23548
rect 13633 23539 13691 23545
rect 8846 23468 8852 23520
rect 8904 23508 8910 23520
rect 9125 23511 9183 23517
rect 9125 23508 9137 23511
rect 8904 23480 9137 23508
rect 8904 23468 8910 23480
rect 9125 23477 9137 23480
rect 9171 23508 9183 23511
rect 9861 23511 9919 23517
rect 9861 23508 9873 23511
rect 9171 23480 9873 23508
rect 9171 23477 9183 23480
rect 9125 23471 9183 23477
rect 9861 23477 9873 23480
rect 9907 23477 9919 23511
rect 9861 23471 9919 23477
rect 10045 23511 10103 23517
rect 10045 23477 10057 23511
rect 10091 23508 10103 23511
rect 10318 23508 10324 23520
rect 10091 23480 10324 23508
rect 10091 23477 10103 23480
rect 10045 23471 10103 23477
rect 10318 23468 10324 23480
rect 10376 23508 10382 23520
rect 13446 23508 13452 23520
rect 10376 23480 13452 23508
rect 10376 23468 10382 23480
rect 13446 23468 13452 23480
rect 13504 23468 13510 23520
rect 14292 23517 14320 23548
rect 17497 23545 17509 23579
rect 17543 23576 17555 23579
rect 17678 23576 17684 23588
rect 17543 23548 17684 23576
rect 17543 23545 17555 23548
rect 17497 23539 17555 23545
rect 17678 23536 17684 23548
rect 17736 23536 17742 23588
rect 20622 23576 20628 23588
rect 20583 23548 20628 23576
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 20824 23576 20852 23616
rect 22066 23616 22192 23644
rect 22066 23576 22094 23616
rect 22186 23604 22192 23616
rect 22244 23644 22250 23656
rect 24489 23647 24547 23653
rect 24489 23644 24501 23647
rect 22244 23616 24501 23644
rect 22244 23604 22250 23616
rect 24489 23613 24501 23616
rect 24535 23613 24547 23647
rect 24489 23607 24547 23613
rect 27982 23604 27988 23656
rect 28040 23644 28046 23656
rect 28261 23647 28319 23653
rect 28261 23644 28273 23647
rect 28040 23616 28273 23644
rect 28040 23604 28046 23616
rect 28261 23613 28273 23616
rect 28307 23613 28319 23647
rect 28261 23607 28319 23613
rect 28721 23647 28779 23653
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 29104 23644 29132 23740
rect 33870 23712 33876 23724
rect 33831 23684 33876 23712
rect 33870 23672 33876 23684
rect 33928 23672 33934 23724
rect 34054 23644 34060 23656
rect 28767 23616 29132 23644
rect 34015 23616 34060 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 34054 23604 34060 23616
rect 34112 23604 34118 23656
rect 30650 23576 30656 23588
rect 20824 23548 22094 23576
rect 25792 23548 30656 23576
rect 14277 23511 14335 23517
rect 14277 23477 14289 23511
rect 14323 23477 14335 23511
rect 14277 23471 14335 23477
rect 16482 23468 16488 23520
rect 16540 23508 16546 23520
rect 18325 23511 18383 23517
rect 18325 23508 18337 23511
rect 16540 23480 18337 23508
rect 16540 23468 16546 23480
rect 18325 23477 18337 23480
rect 18371 23477 18383 23511
rect 18325 23471 18383 23477
rect 22830 23468 22836 23520
rect 22888 23508 22894 23520
rect 22925 23511 22983 23517
rect 22925 23508 22937 23511
rect 22888 23480 22937 23508
rect 22888 23468 22894 23480
rect 22925 23477 22937 23480
rect 22971 23508 22983 23511
rect 25792 23508 25820 23548
rect 30650 23536 30656 23548
rect 30708 23576 30714 23588
rect 30926 23576 30932 23588
rect 30708 23548 30932 23576
rect 30708 23536 30714 23548
rect 30926 23536 30932 23548
rect 30984 23536 30990 23588
rect 22971 23480 25820 23508
rect 25869 23511 25927 23517
rect 22971 23477 22983 23480
rect 22925 23471 22983 23477
rect 25869 23477 25881 23511
rect 25915 23508 25927 23511
rect 26326 23508 26332 23520
rect 25915 23480 26332 23508
rect 25915 23477 25927 23480
rect 25869 23471 25927 23477
rect 26326 23468 26332 23480
rect 26384 23508 26390 23520
rect 27890 23508 27896 23520
rect 26384 23480 27896 23508
rect 26384 23468 26390 23480
rect 27890 23468 27896 23480
rect 27948 23468 27954 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 10134 23304 10140 23316
rect 10095 23276 10140 23304
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 14366 23304 14372 23316
rect 14327 23276 14372 23304
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 15838 23264 15844 23316
rect 15896 23304 15902 23316
rect 16482 23304 16488 23316
rect 15896 23276 16488 23304
rect 15896 23264 15902 23276
rect 16482 23264 16488 23276
rect 16540 23304 16546 23316
rect 17037 23307 17095 23313
rect 17037 23304 17049 23307
rect 16540 23276 17049 23304
rect 16540 23264 16546 23276
rect 17037 23273 17049 23276
rect 17083 23273 17095 23307
rect 17037 23267 17095 23273
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 20349 23307 20407 23313
rect 20349 23304 20361 23307
rect 20128 23276 20361 23304
rect 20128 23264 20134 23276
rect 20349 23273 20361 23276
rect 20395 23273 20407 23307
rect 20349 23267 20407 23273
rect 33873 23307 33931 23313
rect 33873 23273 33885 23307
rect 33919 23304 33931 23307
rect 34054 23304 34060 23316
rect 33919 23276 34060 23304
rect 33919 23273 33931 23276
rect 33873 23267 33931 23273
rect 34054 23264 34060 23276
rect 34112 23264 34118 23316
rect 13722 23196 13728 23248
rect 13780 23236 13786 23248
rect 14274 23236 14280 23248
rect 13780 23208 14280 23236
rect 13780 23196 13786 23208
rect 14274 23196 14280 23208
rect 14332 23196 14338 23248
rect 17221 23239 17279 23245
rect 17221 23205 17233 23239
rect 17267 23205 17279 23239
rect 18414 23236 18420 23248
rect 17221 23199 17279 23205
rect 17328 23208 18420 23236
rect 10318 23168 10324 23180
rect 10060 23140 10324 23168
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 2406 23100 2412 23112
rect 2363 23072 2412 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 2406 23060 2412 23072
rect 2464 23100 2470 23112
rect 2590 23100 2596 23112
rect 2464 23072 2596 23100
rect 2464 23060 2470 23072
rect 2590 23060 2596 23072
rect 2648 23060 2654 23112
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 3694 23100 3700 23112
rect 3007 23072 3700 23100
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 3694 23060 3700 23072
rect 3752 23060 3758 23112
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 9088 23072 9413 23100
rect 9088 23060 9094 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9582 23100 9588 23112
rect 9543 23072 9588 23100
rect 9401 23063 9459 23069
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 10060 23109 10088 23140
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 17126 23168 17132 23180
rect 11808 23140 17132 23168
rect 10045 23103 10103 23109
rect 10045 23069 10057 23103
rect 10091 23069 10103 23103
rect 10045 23063 10103 23069
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 10229 23103 10287 23109
rect 10229 23100 10241 23103
rect 10192 23072 10241 23100
rect 10192 23060 10198 23072
rect 10229 23069 10241 23072
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 10244 23032 10272 23063
rect 10686 23060 10692 23112
rect 10744 23100 10750 23112
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10744 23072 10793 23100
rect 10744 23060 10750 23072
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 10870 23060 10876 23112
rect 10928 23100 10934 23112
rect 11037 23103 11095 23109
rect 11037 23100 11049 23103
rect 10928 23072 11049 23100
rect 10928 23060 10934 23072
rect 11037 23069 11049 23072
rect 11083 23069 11095 23103
rect 11037 23063 11095 23069
rect 11808 23032 11836 23140
rect 17126 23128 17132 23140
rect 17184 23168 17190 23180
rect 17236 23168 17264 23199
rect 17184 23140 17264 23168
rect 17184 23128 17190 23140
rect 12250 23060 12256 23112
rect 12308 23100 12314 23112
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 12308 23072 12725 23100
rect 12308 23060 12314 23072
rect 12713 23069 12725 23072
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23069 12955 23103
rect 12897 23063 12955 23069
rect 12342 23032 12348 23044
rect 10244 23004 11836 23032
rect 12176 23004 12348 23032
rect 2225 22967 2283 22973
rect 2225 22933 2237 22967
rect 2271 22964 2283 22967
rect 3510 22964 3516 22976
rect 2271 22936 3516 22964
rect 2271 22933 2283 22936
rect 2225 22927 2283 22933
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 9493 22967 9551 22973
rect 9493 22933 9505 22967
rect 9539 22964 9551 22967
rect 10042 22964 10048 22976
rect 9539 22936 10048 22964
rect 9539 22933 9551 22936
rect 9493 22927 9551 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 12176 22973 12204 23004
rect 12342 22992 12348 23004
rect 12400 23032 12406 23044
rect 12912 23032 12940 23063
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 14277 23103 14335 23109
rect 14277 23100 14289 23103
rect 13872 23072 14289 23100
rect 13872 23060 13878 23072
rect 14277 23069 14289 23072
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 16114 23060 16120 23112
rect 16172 23100 16178 23112
rect 16209 23103 16267 23109
rect 16209 23100 16221 23103
rect 16172 23072 16221 23100
rect 16172 23060 16178 23072
rect 16209 23069 16221 23072
rect 16255 23069 16267 23103
rect 17328 23100 17356 23208
rect 18414 23196 18420 23208
rect 18472 23196 18478 23248
rect 20162 23236 20168 23248
rect 20123 23208 20168 23236
rect 20162 23196 20168 23208
rect 20220 23196 20226 23248
rect 22094 23236 22100 23248
rect 20272 23208 22100 23236
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 20272 23168 20300 23208
rect 22094 23196 22100 23208
rect 22152 23196 22158 23248
rect 26786 23236 26792 23248
rect 26747 23208 26792 23236
rect 26786 23196 26792 23208
rect 26844 23196 26850 23248
rect 31021 23239 31079 23245
rect 31021 23205 31033 23239
rect 31067 23236 31079 23239
rect 31067 23208 31800 23236
rect 31067 23205 31079 23208
rect 31021 23199 31079 23205
rect 18187 23140 20300 23168
rect 20441 23171 20499 23177
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 20441 23137 20453 23171
rect 20487 23168 20499 23171
rect 21082 23168 21088 23180
rect 20487 23140 21088 23168
rect 20487 23137 20499 23140
rect 20441 23131 20499 23137
rect 21082 23128 21088 23140
rect 21140 23128 21146 23180
rect 22278 23168 22284 23180
rect 21468 23140 22284 23168
rect 17770 23100 17776 23112
rect 16209 23063 16267 23069
rect 16316 23072 17356 23100
rect 17731 23072 17776 23100
rect 16316 23032 16344 23072
rect 17770 23060 17776 23072
rect 17828 23060 17834 23112
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23100 18015 23103
rect 18046 23100 18052 23112
rect 18003 23072 18052 23100
rect 18003 23069 18015 23072
rect 17957 23063 18015 23069
rect 18046 23060 18052 23072
rect 18104 23060 18110 23112
rect 21468 23109 21496 23140
rect 20533 23103 20591 23109
rect 20533 23069 20545 23103
rect 20579 23069 20591 23103
rect 20533 23063 20591 23069
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 12400 23004 16344 23032
rect 16393 23035 16451 23041
rect 12400 22992 12406 23004
rect 16393 23001 16405 23035
rect 16439 23032 16451 23035
rect 16853 23035 16911 23041
rect 16853 23032 16865 23035
rect 16439 23004 16865 23032
rect 16439 23001 16451 23004
rect 16393 22995 16451 23001
rect 16853 23001 16865 23004
rect 16899 23032 16911 23035
rect 17862 23032 17868 23044
rect 16899 23004 17868 23032
rect 16899 23001 16911 23004
rect 16853 22995 16911 23001
rect 17862 22992 17868 23004
rect 17920 22992 17926 23044
rect 18693 23035 18751 23041
rect 18693 23001 18705 23035
rect 18739 23001 18751 23035
rect 18693 22995 18751 23001
rect 12161 22967 12219 22973
rect 12161 22933 12173 22967
rect 12207 22933 12219 22967
rect 12161 22927 12219 22933
rect 12897 22967 12955 22973
rect 12897 22933 12909 22967
rect 12943 22964 12955 22967
rect 14734 22964 14740 22976
rect 12943 22936 14740 22964
rect 12943 22933 12955 22936
rect 12897 22927 12955 22933
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 17034 22924 17040 22976
rect 17092 22973 17098 22976
rect 17092 22967 17111 22973
rect 17099 22964 17111 22967
rect 17678 22964 17684 22976
rect 17099 22936 17684 22964
rect 17099 22933 17111 22936
rect 17092 22927 17111 22933
rect 17092 22924 17098 22927
rect 17678 22924 17684 22936
rect 17736 22964 17742 22976
rect 18708 22964 18736 22995
rect 20346 22992 20352 23044
rect 20404 23032 20410 23044
rect 20548 23032 20576 23063
rect 20404 23004 20576 23032
rect 21836 23032 21864 23140
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 23566 23168 23572 23180
rect 23479 23140 23572 23168
rect 23492 23109 23520 23140
rect 23566 23128 23572 23140
rect 23624 23168 23630 23180
rect 24854 23168 24860 23180
rect 23624 23140 24860 23168
rect 23624 23128 23630 23140
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 26326 23168 26332 23180
rect 26287 23140 26332 23168
rect 26326 23128 26332 23140
rect 26384 23128 26390 23180
rect 30374 23128 30380 23180
rect 30432 23168 30438 23180
rect 31772 23177 31800 23208
rect 30561 23171 30619 23177
rect 30561 23168 30573 23171
rect 30432 23140 30573 23168
rect 30432 23128 30438 23140
rect 30561 23137 30573 23140
rect 30607 23137 30619 23171
rect 30561 23131 30619 23137
rect 31757 23171 31815 23177
rect 31757 23137 31769 23171
rect 31803 23137 31815 23171
rect 31757 23131 31815 23137
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23100 21971 23103
rect 22925 23103 22983 23109
rect 22925 23100 22937 23103
rect 21959 23072 22937 23100
rect 21959 23069 21971 23072
rect 21913 23063 21971 23069
rect 22925 23069 22937 23072
rect 22971 23069 22983 23103
rect 22925 23063 22983 23069
rect 23477 23103 23535 23109
rect 23477 23069 23489 23103
rect 23523 23069 23535 23103
rect 23658 23100 23664 23112
rect 23619 23072 23664 23100
rect 23477 23063 23535 23069
rect 23658 23060 23664 23072
rect 23716 23100 23722 23112
rect 24302 23100 24308 23112
rect 23716 23072 24308 23100
rect 23716 23060 23722 23072
rect 24302 23060 24308 23072
rect 24360 23060 24366 23112
rect 26421 23103 26479 23109
rect 26421 23069 26433 23103
rect 26467 23100 26479 23103
rect 26970 23100 26976 23112
rect 26467 23072 26976 23100
rect 26467 23069 26479 23072
rect 26421 23063 26479 23069
rect 26970 23060 26976 23072
rect 27028 23100 27034 23112
rect 30653 23103 30711 23109
rect 30653 23100 30665 23103
rect 27028 23072 30665 23100
rect 27028 23060 27034 23072
rect 30653 23069 30665 23072
rect 30699 23100 30711 23103
rect 30742 23100 30748 23112
rect 30699 23072 30748 23100
rect 30699 23069 30711 23072
rect 30653 23063 30711 23069
rect 30742 23060 30748 23072
rect 30800 23060 30806 23112
rect 31846 23100 31852 23112
rect 31807 23072 31852 23100
rect 31846 23060 31852 23072
rect 31904 23060 31910 23112
rect 33781 23103 33839 23109
rect 33781 23069 33793 23103
rect 33827 23100 33839 23103
rect 33870 23100 33876 23112
rect 33827 23072 33876 23100
rect 33827 23069 33839 23072
rect 33781 23063 33839 23069
rect 33870 23060 33876 23072
rect 33928 23060 33934 23112
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23100 37887 23103
rect 38286 23100 38292 23112
rect 37875 23072 38292 23100
rect 37875 23069 37887 23072
rect 37829 23063 37887 23069
rect 38286 23060 38292 23072
rect 38344 23060 38350 23112
rect 22097 23035 22155 23041
rect 22097 23032 22109 23035
rect 21836 23004 22109 23032
rect 20404 22992 20410 23004
rect 22097 23001 22109 23004
rect 22143 23001 22155 23035
rect 22097 22995 22155 23001
rect 22281 23035 22339 23041
rect 22281 23001 22293 23035
rect 22327 23032 22339 23035
rect 24210 23032 24216 23044
rect 22327 23004 24216 23032
rect 22327 23001 22339 23004
rect 22281 22995 22339 23001
rect 24210 22992 24216 23004
rect 24268 22992 24274 23044
rect 17736 22936 18736 22964
rect 17736 22924 17742 22936
rect 18782 22924 18788 22976
rect 18840 22964 18846 22976
rect 21269 22967 21327 22973
rect 18840 22936 18885 22964
rect 18840 22924 18846 22936
rect 21269 22933 21281 22967
rect 21315 22964 21327 22967
rect 21910 22964 21916 22976
rect 21315 22936 21916 22964
rect 21315 22933 21327 22936
rect 21269 22927 21327 22933
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 22738 22964 22744 22976
rect 22699 22936 22744 22964
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 23661 22967 23719 22973
rect 23661 22933 23673 22967
rect 23707 22964 23719 22967
rect 23750 22964 23756 22976
rect 23707 22936 23756 22964
rect 23707 22933 23719 22936
rect 23661 22927 23719 22933
rect 23750 22924 23756 22936
rect 23808 22924 23814 22976
rect 31018 22924 31024 22976
rect 31076 22964 31082 22976
rect 31481 22967 31539 22973
rect 31481 22964 31493 22967
rect 31076 22936 31493 22964
rect 31076 22924 31082 22936
rect 31481 22933 31493 22936
rect 31527 22933 31539 22967
rect 31481 22927 31539 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 12621 22763 12679 22769
rect 12621 22760 12633 22763
rect 8956 22732 12633 22760
rect 3510 22692 3516 22704
rect 3471 22664 3516 22692
rect 3510 22652 3516 22664
rect 3568 22652 3574 22704
rect 3694 22584 3700 22636
rect 3752 22624 3758 22636
rect 8956 22633 8984 22732
rect 12621 22729 12633 22732
rect 12667 22760 12679 22763
rect 13722 22760 13728 22772
rect 12667 22732 13728 22760
rect 12667 22729 12679 22732
rect 12621 22723 12679 22729
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 15470 22760 15476 22772
rect 15431 22732 15476 22760
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 17770 22760 17776 22772
rect 17267 22732 17776 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 18230 22760 18236 22772
rect 18191 22732 18236 22760
rect 18230 22720 18236 22732
rect 18288 22720 18294 22772
rect 18417 22763 18475 22769
rect 18417 22729 18429 22763
rect 18463 22729 18475 22763
rect 18417 22723 18475 22729
rect 15105 22695 15163 22701
rect 15105 22661 15117 22695
rect 15151 22692 15163 22695
rect 16114 22692 16120 22704
rect 15151 22664 16120 22692
rect 15151 22661 15163 22664
rect 15105 22655 15163 22661
rect 8941 22627 8999 22633
rect 3752 22596 3797 22624
rect 3752 22584 3758 22596
rect 8941 22593 8953 22627
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 12805 22627 12863 22633
rect 12805 22624 12817 22627
rect 12492 22596 12817 22624
rect 12492 22584 12498 22596
rect 12805 22593 12817 22596
rect 12851 22593 12863 22627
rect 12805 22587 12863 22593
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 14826 22624 14832 22636
rect 13504 22596 14832 22624
rect 13504 22584 13510 22596
rect 14826 22584 14832 22596
rect 14884 22584 14890 22636
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 1854 22556 1860 22568
rect 1815 22528 1860 22556
rect 1854 22516 1860 22528
rect 1912 22516 1918 22568
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 9309 22559 9367 22565
rect 9309 22525 9321 22559
rect 9355 22556 9367 22559
rect 9582 22556 9588 22568
rect 9355 22528 9588 22556
rect 9355 22525 9367 22528
rect 9309 22519 9367 22525
rect 9048 22488 9076 22519
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 15304 22556 15332 22587
rect 15654 22584 15660 22636
rect 15712 22624 15718 22636
rect 16040 22633 16068 22664
rect 16114 22652 16120 22664
rect 16172 22652 16178 22704
rect 17586 22652 17592 22704
rect 17644 22692 17650 22704
rect 17862 22692 17868 22704
rect 17644 22664 17868 22692
rect 17644 22652 17650 22664
rect 17862 22652 17868 22664
rect 17920 22692 17926 22704
rect 18432 22692 18460 22723
rect 21910 22720 21916 22772
rect 21968 22760 21974 22772
rect 30558 22760 30564 22772
rect 21968 22732 23428 22760
rect 30519 22732 30564 22760
rect 21968 22720 21974 22732
rect 22278 22692 22284 22704
rect 17920 22664 18460 22692
rect 18524 22664 22284 22692
rect 17920 22652 17926 22664
rect 15921 22627 15979 22633
rect 15921 22624 15933 22627
rect 15712 22596 15933 22624
rect 15712 22584 15718 22596
rect 15921 22593 15933 22596
rect 15967 22593 15979 22627
rect 15921 22587 15979 22593
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22624 16083 22627
rect 16850 22624 16856 22636
rect 16071 22596 16105 22624
rect 16811 22596 16856 22624
rect 16071 22593 16083 22596
rect 16025 22587 16083 22593
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 17402 22624 17408 22636
rect 17083 22596 17408 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 18358 22627 18416 22633
rect 18358 22624 18370 22627
rect 17512 22596 18370 22624
rect 12768 22528 15332 22556
rect 12768 22516 12774 22528
rect 9858 22488 9864 22500
rect 9048 22460 9864 22488
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 15304 22488 15332 22528
rect 17512 22488 17540 22596
rect 18358 22593 18370 22596
rect 18404 22624 18416 22627
rect 18524 22624 18552 22664
rect 22278 22652 22284 22664
rect 22336 22652 22342 22704
rect 22456 22695 22514 22701
rect 22456 22661 22468 22695
rect 22502 22692 22514 22695
rect 22738 22692 22744 22704
rect 22502 22664 22744 22692
rect 22502 22661 22514 22664
rect 22456 22655 22514 22661
rect 22738 22652 22744 22664
rect 22796 22652 22802 22704
rect 18404 22596 18552 22624
rect 20441 22627 20499 22633
rect 18404 22593 18416 22596
rect 18358 22587 18416 22593
rect 20441 22593 20453 22627
rect 20487 22593 20499 22627
rect 20441 22587 20499 22593
rect 18877 22559 18935 22565
rect 18877 22525 18889 22559
rect 18923 22556 18935 22559
rect 19978 22556 19984 22568
rect 18923 22528 19984 22556
rect 18923 22525 18935 22528
rect 18877 22519 18935 22525
rect 19978 22516 19984 22528
rect 20036 22516 20042 22568
rect 20456 22556 20484 22587
rect 20530 22584 20536 22636
rect 20588 22624 20594 22636
rect 20588 22596 20633 22624
rect 20588 22584 20594 22596
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 22186 22624 22192 22636
rect 20772 22596 21496 22624
rect 22147 22596 22192 22624
rect 20772 22584 20778 22596
rect 21358 22556 21364 22568
rect 20456 22528 21364 22556
rect 21358 22516 21364 22528
rect 21416 22516 21422 22568
rect 21468 22556 21496 22596
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 23400 22624 23428 22732
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 24762 22692 24768 22704
rect 24723 22664 24768 22692
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 29546 22624 29552 22636
rect 22296 22596 23244 22624
rect 23400 22596 29552 22624
rect 22296 22556 22324 22596
rect 21468 22528 22324 22556
rect 23216 22556 23244 22596
rect 29546 22584 29552 22596
rect 29604 22584 29610 22636
rect 30374 22584 30380 22636
rect 30432 22624 30438 22636
rect 30502 22627 30560 22633
rect 30502 22624 30514 22627
rect 30432 22596 30514 22624
rect 30432 22584 30438 22596
rect 30502 22593 30514 22596
rect 30548 22593 30560 22627
rect 31018 22624 31024 22636
rect 30979 22596 31024 22624
rect 30502 22587 30560 22593
rect 31018 22584 31024 22596
rect 31076 22584 31082 22636
rect 37458 22624 37464 22636
rect 37419 22596 37464 22624
rect 37458 22584 37464 22596
rect 37516 22624 37522 22636
rect 37734 22624 37740 22636
rect 37516 22596 37740 22624
rect 37516 22584 37522 22596
rect 37734 22584 37740 22596
rect 37792 22584 37798 22636
rect 29270 22556 29276 22568
rect 23216 22528 29276 22556
rect 29270 22516 29276 22528
rect 29328 22516 29334 22568
rect 30650 22516 30656 22568
rect 30708 22556 30714 22568
rect 30929 22559 30987 22565
rect 30929 22556 30941 22559
rect 30708 22528 30941 22556
rect 30708 22516 30714 22528
rect 30929 22525 30941 22528
rect 30975 22525 30987 22559
rect 30929 22519 30987 22525
rect 23566 22488 23572 22500
rect 15304 22460 17540 22488
rect 23479 22460 23572 22488
rect 23566 22448 23572 22460
rect 23624 22488 23630 22500
rect 24762 22488 24768 22500
rect 23624 22460 24768 22488
rect 23624 22448 23630 22460
rect 24762 22448 24768 22460
rect 24820 22448 24826 22500
rect 24949 22491 25007 22497
rect 24949 22457 24961 22491
rect 24995 22488 25007 22491
rect 25866 22488 25872 22500
rect 24995 22460 25872 22488
rect 24995 22457 25007 22460
rect 24949 22451 25007 22457
rect 25866 22448 25872 22460
rect 25924 22448 25930 22500
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 15933 22423 15991 22429
rect 15933 22420 15945 22423
rect 15896 22392 15945 22420
rect 15896 22380 15902 22392
rect 15933 22389 15945 22392
rect 15979 22389 15991 22423
rect 15933 22383 15991 22389
rect 16301 22423 16359 22429
rect 16301 22389 16313 22423
rect 16347 22420 16359 22423
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 16347 22392 16865 22420
rect 16347 22389 16359 22392
rect 16301 22383 16359 22389
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 16853 22383 16911 22389
rect 18414 22380 18420 22432
rect 18472 22420 18478 22432
rect 18785 22423 18843 22429
rect 18785 22420 18797 22423
rect 18472 22392 18797 22420
rect 18472 22380 18478 22392
rect 18785 22389 18797 22392
rect 18831 22389 18843 22423
rect 18785 22383 18843 22389
rect 20901 22423 20959 22429
rect 20901 22389 20913 22423
rect 20947 22420 20959 22423
rect 23382 22420 23388 22432
rect 20947 22392 23388 22420
rect 20947 22389 20959 22392
rect 20901 22383 20959 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 30374 22420 30380 22432
rect 30335 22392 30380 22420
rect 30374 22380 30380 22392
rect 30432 22380 30438 22432
rect 37553 22423 37611 22429
rect 37553 22389 37565 22423
rect 37599 22420 37611 22423
rect 38102 22420 38108 22432
rect 37599 22392 38108 22420
rect 37599 22389 37611 22392
rect 37553 22383 37611 22389
rect 38102 22380 38108 22392
rect 38160 22380 38166 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 13078 22176 13084 22228
rect 13136 22216 13142 22228
rect 13357 22219 13415 22225
rect 13357 22216 13369 22219
rect 13136 22188 13369 22216
rect 13136 22176 13142 22188
rect 13357 22185 13369 22188
rect 13403 22185 13415 22219
rect 13357 22179 13415 22185
rect 13725 22219 13783 22225
rect 13725 22185 13737 22219
rect 13771 22216 13783 22219
rect 14090 22216 14096 22228
rect 13771 22188 14096 22216
rect 13771 22185 13783 22188
rect 13725 22179 13783 22185
rect 14090 22176 14096 22188
rect 14148 22216 14154 22228
rect 14921 22219 14979 22225
rect 14921 22216 14933 22219
rect 14148 22188 14933 22216
rect 14148 22176 14154 22188
rect 14921 22185 14933 22188
rect 14967 22216 14979 22219
rect 15010 22216 15016 22228
rect 14967 22188 15016 22216
rect 14967 22185 14979 22188
rect 14921 22179 14979 22185
rect 15010 22176 15016 22188
rect 15068 22176 15074 22228
rect 15470 22176 15476 22228
rect 15528 22216 15534 22228
rect 15565 22219 15623 22225
rect 15565 22216 15577 22219
rect 15528 22188 15577 22216
rect 15528 22176 15534 22188
rect 15565 22185 15577 22188
rect 15611 22185 15623 22219
rect 15565 22179 15623 22185
rect 20165 22219 20223 22225
rect 20165 22185 20177 22219
rect 20211 22216 20223 22219
rect 20530 22216 20536 22228
rect 20211 22188 20536 22216
rect 20211 22185 20223 22188
rect 20165 22179 20223 22185
rect 20530 22176 20536 22188
rect 20588 22176 20594 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 20809 22219 20867 22225
rect 20809 22216 20821 22219
rect 20772 22188 20821 22216
rect 20772 22176 20778 22188
rect 20809 22185 20821 22188
rect 20855 22216 20867 22219
rect 21174 22216 21180 22228
rect 20855 22188 21180 22216
rect 20855 22185 20867 22188
rect 20809 22179 20867 22185
rect 21174 22176 21180 22188
rect 21232 22176 21238 22228
rect 26050 22176 26056 22228
rect 26108 22216 26114 22228
rect 28626 22216 28632 22228
rect 26108 22188 28632 22216
rect 26108 22176 26114 22188
rect 28626 22176 28632 22188
rect 28684 22176 28690 22228
rect 30466 22176 30472 22228
rect 30524 22216 30530 22228
rect 31113 22219 31171 22225
rect 31113 22216 31125 22219
rect 30524 22188 31125 22216
rect 30524 22176 30530 22188
rect 31113 22185 31125 22188
rect 31159 22185 31171 22219
rect 31113 22179 31171 22185
rect 27172 22120 27568 22148
rect 2774 22040 2780 22092
rect 2832 22080 2838 22092
rect 2832 22052 2877 22080
rect 2832 22040 2838 22052
rect 8662 22040 8668 22092
rect 8720 22080 8726 22092
rect 12805 22083 12863 22089
rect 12805 22080 12817 22083
rect 8720 22052 10824 22080
rect 8720 22040 8726 22052
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 10686 22012 10692 22024
rect 10647 21984 10692 22012
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 10796 22012 10824 22052
rect 12406 22052 12817 22080
rect 12406 22012 12434 22052
rect 12805 22049 12817 22052
rect 12851 22080 12863 22083
rect 14182 22080 14188 22092
rect 12851 22052 14188 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 14734 22080 14740 22092
rect 14695 22052 14740 22080
rect 14734 22040 14740 22052
rect 14792 22080 14798 22092
rect 15654 22080 15660 22092
rect 14792 22052 15660 22080
rect 14792 22040 14798 22052
rect 15654 22040 15660 22052
rect 15712 22040 15718 22092
rect 17402 22080 17408 22092
rect 17363 22052 17408 22080
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 17862 22080 17868 22092
rect 17823 22052 17868 22080
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 24210 22040 24216 22092
rect 24268 22080 24274 22092
rect 24268 22052 24992 22080
rect 24268 22040 24274 22052
rect 10796 21984 12434 22012
rect 12710 21972 12716 22024
rect 12768 21972 12774 22024
rect 13170 21972 13176 22024
rect 13228 22012 13234 22024
rect 13357 22015 13415 22021
rect 13357 22012 13369 22015
rect 13228 21984 13369 22012
rect 13228 21972 13234 21984
rect 13357 21981 13369 21984
rect 13403 21981 13415 22015
rect 13357 21975 13415 21981
rect 13446 21972 13452 22024
rect 13504 22012 13510 22024
rect 14918 22012 14924 22024
rect 13504 21984 13549 22012
rect 14879 21984 14924 22012
rect 13504 21972 13510 21984
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 15010 21972 15016 22024
rect 15068 22012 15074 22024
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 15068 21984 15853 22012
rect 15068 21972 15074 21984
rect 15841 21981 15853 21984
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 17313 22015 17371 22021
rect 17313 21981 17325 22015
rect 17359 21981 17371 22015
rect 20070 22012 20076 22024
rect 20031 21984 20076 22012
rect 17313 21975 17371 21981
rect 1765 21947 1823 21953
rect 1765 21913 1777 21947
rect 1811 21944 1823 21947
rect 2406 21944 2412 21956
rect 1811 21916 2412 21944
rect 1811 21913 1823 21916
rect 1765 21907 1823 21913
rect 2406 21904 2412 21916
rect 2464 21904 2470 21956
rect 10042 21904 10048 21956
rect 10100 21944 10106 21956
rect 10934 21947 10992 21953
rect 10934 21944 10946 21947
rect 10100 21916 10946 21944
rect 10100 21904 10106 21916
rect 10934 21913 10946 21916
rect 10980 21913 10992 21947
rect 10934 21907 10992 21913
rect 12621 21947 12679 21953
rect 12621 21913 12633 21947
rect 12667 21944 12679 21947
rect 12728 21944 12756 21972
rect 12986 21944 12992 21956
rect 12667 21916 12992 21944
rect 12667 21913 12679 21916
rect 12621 21907 12679 21913
rect 12986 21904 12992 21916
rect 13044 21904 13050 21956
rect 14366 21904 14372 21956
rect 14424 21944 14430 21956
rect 14461 21947 14519 21953
rect 14461 21944 14473 21947
rect 14424 21916 14473 21944
rect 14424 21904 14430 21916
rect 14461 21913 14473 21916
rect 14507 21913 14519 21947
rect 15562 21944 15568 21956
rect 15523 21916 15568 21944
rect 14461 21907 14519 21913
rect 15562 21904 15568 21916
rect 15620 21904 15626 21956
rect 12069 21879 12127 21885
rect 12069 21845 12081 21879
rect 12115 21876 12127 21879
rect 12434 21876 12440 21888
rect 12115 21848 12440 21876
rect 12115 21845 12127 21848
rect 12069 21839 12127 21845
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 15102 21876 15108 21888
rect 15063 21848 15108 21876
rect 15102 21836 15108 21848
rect 15160 21836 15166 21888
rect 16025 21879 16083 21885
rect 16025 21845 16037 21879
rect 16071 21876 16083 21879
rect 17328 21876 17356 21975
rect 20070 21972 20076 21984
rect 20128 21972 20134 22024
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 22012 20315 22015
rect 20898 22012 20904 22024
rect 20303 21984 20904 22012
rect 20303 21981 20315 21984
rect 20257 21975 20315 21981
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21085 22015 21143 22021
rect 21085 21981 21097 22015
rect 21131 22012 21143 22015
rect 21266 22012 21272 22024
rect 21131 21984 21272 22012
rect 21131 21981 21143 21984
rect 21085 21975 21143 21981
rect 21266 21972 21272 21984
rect 21324 21972 21330 22024
rect 23661 22015 23719 22021
rect 23661 21981 23673 22015
rect 23707 22012 23719 22015
rect 23750 22012 23756 22024
rect 23707 21984 23756 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 23750 21972 23756 21984
rect 23808 21972 23814 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 24854 22012 24860 22024
rect 24815 21984 24860 22012
rect 23845 21975 23903 21981
rect 18506 21904 18512 21956
rect 18564 21944 18570 21956
rect 23860 21944 23888 21975
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 24964 22012 24992 22052
rect 25866 22040 25872 22092
rect 25924 22080 25930 22092
rect 27172 22080 27200 22120
rect 27338 22080 27344 22092
rect 25924 22052 27200 22080
rect 27299 22052 27344 22080
rect 25924 22040 25930 22052
rect 27338 22040 27344 22052
rect 27396 22040 27402 22092
rect 26881 22015 26939 22021
rect 26881 22012 26893 22015
rect 24964 21984 26893 22012
rect 26881 21981 26893 21984
rect 26927 21981 26939 22015
rect 26881 21975 26939 21981
rect 27065 22015 27123 22021
rect 27065 21981 27077 22015
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 24118 21944 24124 21956
rect 18564 21916 24124 21944
rect 18564 21904 18570 21916
rect 24118 21904 24124 21916
rect 24176 21904 24182 21956
rect 24394 21904 24400 21956
rect 24452 21944 24458 21956
rect 25102 21947 25160 21953
rect 25102 21944 25114 21947
rect 24452 21916 25114 21944
rect 24452 21904 24458 21916
rect 25102 21913 25114 21916
rect 25148 21913 25160 21947
rect 25102 21907 25160 21913
rect 16071 21848 17356 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 17681 21879 17739 21885
rect 17681 21876 17693 21879
rect 17552 21848 17693 21876
rect 17552 21836 17558 21848
rect 17681 21845 17693 21848
rect 17727 21876 17739 21879
rect 23658 21876 23664 21888
rect 17727 21848 23664 21876
rect 17727 21845 17739 21848
rect 17681 21839 17739 21845
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 23845 21879 23903 21885
rect 23845 21845 23857 21879
rect 23891 21876 23903 21879
rect 23934 21876 23940 21888
rect 23891 21848 23940 21876
rect 23891 21845 23903 21848
rect 23845 21839 23903 21845
rect 23934 21836 23940 21848
rect 23992 21836 23998 21888
rect 26234 21876 26240 21888
rect 26195 21848 26240 21876
rect 26234 21836 26240 21848
rect 26292 21836 26298 21888
rect 27080 21876 27108 21975
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 27433 22015 27491 22021
rect 27212 21984 27257 22012
rect 27212 21972 27218 21984
rect 27433 21981 27445 22015
rect 27479 22012 27491 22015
rect 27540 22012 27568 22120
rect 37182 22080 37188 22092
rect 37143 22052 37188 22080
rect 37182 22040 37188 22052
rect 37240 22040 37246 22092
rect 38102 22080 38108 22092
rect 38063 22052 38108 22080
rect 38102 22040 38108 22052
rect 38160 22040 38166 22092
rect 38286 22080 38292 22092
rect 38247 22052 38292 22080
rect 38286 22040 38292 22052
rect 38344 22040 38350 22092
rect 27479 21984 27568 22012
rect 27479 21981 27491 21984
rect 27433 21975 27491 21981
rect 27706 21972 27712 22024
rect 27764 22012 27770 22024
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 27764 21984 29745 22012
rect 27764 21972 27770 21984
rect 29733 21981 29745 21984
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 29638 21904 29644 21956
rect 29696 21944 29702 21956
rect 29978 21947 30036 21953
rect 29978 21944 29990 21947
rect 29696 21916 29990 21944
rect 29696 21904 29702 21916
rect 29978 21913 29990 21916
rect 30024 21913 30036 21947
rect 29978 21907 30036 21913
rect 27798 21876 27804 21888
rect 27080 21848 27804 21876
rect 27798 21836 27804 21848
rect 27856 21836 27862 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2406 21672 2412 21684
rect 2367 21644 2412 21672
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 14001 21675 14059 21681
rect 14001 21641 14013 21675
rect 14047 21672 14059 21675
rect 15105 21675 15163 21681
rect 14047 21644 15056 21672
rect 14047 21641 14059 21644
rect 14001 21635 14059 21641
rect 9033 21607 9091 21613
rect 9033 21573 9045 21607
rect 9079 21604 9091 21607
rect 12069 21607 12127 21613
rect 9079 21576 9720 21604
rect 9079 21573 9091 21576
rect 9033 21567 9091 21573
rect 1578 21496 1584 21548
rect 1636 21536 1642 21548
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 1636 21508 1685 21536
rect 1636 21496 1642 21508
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 2682 21536 2688 21548
rect 2547 21508 2688 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 2682 21496 2688 21508
rect 2740 21496 2746 21548
rect 2774 21496 2780 21548
rect 2832 21536 2838 21548
rect 2961 21539 3019 21545
rect 2961 21536 2973 21539
rect 2832 21508 2973 21536
rect 2832 21496 2838 21508
rect 2961 21505 2973 21508
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 8757 21539 8815 21545
rect 8757 21536 8769 21539
rect 8720 21508 8769 21536
rect 8720 21496 8726 21508
rect 8757 21505 8769 21508
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 8846 21496 8852 21548
rect 8904 21536 8910 21548
rect 8904 21508 8949 21536
rect 8904 21496 8910 21508
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9692 21545 9720 21576
rect 12069 21573 12081 21607
rect 12115 21604 12127 21607
rect 12434 21604 12440 21616
rect 12115 21576 12440 21604
rect 12115 21573 12127 21576
rect 12069 21567 12127 21573
rect 12434 21564 12440 21576
rect 12492 21604 12498 21616
rect 12713 21607 12771 21613
rect 12713 21604 12725 21607
rect 12492 21576 12725 21604
rect 12492 21564 12498 21576
rect 12713 21573 12725 21576
rect 12759 21604 12771 21607
rect 15028 21604 15056 21644
rect 15105 21641 15117 21675
rect 15151 21672 15163 21675
rect 15562 21672 15568 21684
rect 15151 21644 15568 21672
rect 15151 21641 15163 21644
rect 15105 21635 15163 21641
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 17144 21644 19932 21672
rect 17144 21604 17172 21644
rect 12759 21576 14412 21604
rect 15028 21576 17172 21604
rect 12759 21573 12771 21576
rect 12713 21567 12771 21573
rect 14384 21548 14412 21576
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 17313 21607 17371 21613
rect 17313 21604 17325 21607
rect 17276 21576 17325 21604
rect 17276 21564 17282 21576
rect 17313 21573 17325 21576
rect 17359 21573 17371 21607
rect 17313 21567 17371 21573
rect 17497 21607 17555 21613
rect 17497 21573 17509 21607
rect 17543 21604 17555 21607
rect 17954 21604 17960 21616
rect 17543 21576 17960 21604
rect 17543 21573 17555 21576
rect 17497 21567 17555 21573
rect 9493 21539 9551 21545
rect 9493 21536 9505 21539
rect 9180 21508 9505 21536
rect 9180 21496 9186 21508
rect 9493 21505 9505 21508
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21505 9735 21539
rect 9677 21499 9735 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 11974 21536 11980 21548
rect 11931 21508 11980 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 11974 21496 11980 21508
rect 12032 21536 12038 21548
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 12032 21508 13185 21536
rect 12032 21496 12038 21508
rect 13173 21505 13185 21508
rect 13219 21505 13231 21539
rect 13173 21499 13231 21505
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 13909 21539 13967 21545
rect 13909 21536 13921 21539
rect 13872 21508 13921 21536
rect 13872 21496 13878 21508
rect 13909 21505 13921 21508
rect 13955 21505 13967 21539
rect 14090 21536 14096 21548
rect 14051 21508 14096 21536
rect 13909 21499 13967 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 14424 21508 14565 21536
rect 14424 21496 14430 21508
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 15102 21496 15108 21548
rect 15160 21536 15166 21548
rect 15565 21539 15623 21545
rect 15565 21536 15577 21539
rect 15160 21508 15577 21536
rect 15160 21496 15166 21508
rect 15565 21505 15577 21508
rect 15611 21505 15623 21539
rect 15565 21499 15623 21505
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21536 15899 21539
rect 15930 21536 15936 21548
rect 15887 21508 15936 21536
rect 15887 21505 15899 21508
rect 15841 21499 15899 21505
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 17512 21536 17540 21567
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 17328 21508 17540 21536
rect 18785 21539 18843 21545
rect 2700 21468 2728 21496
rect 3602 21468 3608 21480
rect 2700 21440 3608 21468
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 9033 21471 9091 21477
rect 9033 21437 9045 21471
rect 9079 21468 9091 21471
rect 9582 21468 9588 21480
rect 9079 21440 9588 21468
rect 9079 21437 9091 21440
rect 9033 21431 9091 21437
rect 9582 21428 9588 21440
rect 9640 21428 9646 21480
rect 12986 21468 12992 21480
rect 12947 21440 12992 21468
rect 12986 21428 12992 21440
rect 13044 21428 13050 21480
rect 14458 21428 14464 21480
rect 14516 21468 14522 21480
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 14516 21440 14841 21468
rect 14516 21428 14522 21440
rect 14829 21437 14841 21440
rect 14875 21468 14887 21471
rect 14918 21468 14924 21480
rect 14875 21440 14924 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 15528 21440 15669 21468
rect 15528 21428 15534 21440
rect 15657 21437 15669 21440
rect 15703 21437 15715 21471
rect 15657 21431 15715 21437
rect 13814 21400 13820 21412
rect 12360 21372 13820 21400
rect 12360 21344 12388 21372
rect 13814 21360 13820 21372
rect 13872 21360 13878 21412
rect 14182 21360 14188 21412
rect 14240 21400 14246 21412
rect 15194 21400 15200 21412
rect 14240 21372 15200 21400
rect 14240 21360 14246 21372
rect 15194 21360 15200 21372
rect 15252 21360 15258 21412
rect 15565 21403 15623 21409
rect 15565 21369 15577 21403
rect 15611 21400 15623 21403
rect 17328 21400 17356 21508
rect 18785 21505 18797 21539
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21536 19027 21539
rect 19794 21536 19800 21548
rect 19015 21508 19800 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 18800 21468 18828 21499
rect 19794 21496 19800 21508
rect 19852 21496 19858 21548
rect 19904 21536 19932 21644
rect 20898 21632 20904 21684
rect 20956 21672 20962 21684
rect 20993 21675 21051 21681
rect 20993 21672 21005 21675
rect 20956 21644 21005 21672
rect 20956 21632 20962 21644
rect 20993 21641 21005 21644
rect 21039 21641 21051 21675
rect 21358 21672 21364 21684
rect 21319 21644 21364 21672
rect 20993 21635 21051 21641
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 24026 21632 24032 21684
rect 24084 21672 24090 21684
rect 24394 21672 24400 21684
rect 24084 21644 24256 21672
rect 24355 21644 24400 21672
rect 24084 21632 24090 21644
rect 23198 21564 23204 21616
rect 23256 21604 23262 21616
rect 24228 21604 24256 21644
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 24854 21632 24860 21684
rect 24912 21672 24918 21684
rect 27706 21672 27712 21684
rect 24912 21644 27712 21672
rect 24912 21632 24918 21644
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 29638 21672 29644 21684
rect 29599 21644 29644 21672
rect 29638 21632 29644 21644
rect 29696 21632 29702 21684
rect 27154 21604 27160 21616
rect 23256 21576 24072 21604
rect 24228 21576 27160 21604
rect 23256 21564 23262 21576
rect 20346 21536 20352 21548
rect 19904 21508 20352 21536
rect 20346 21496 20352 21508
rect 20404 21536 20410 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20404 21508 20913 21536
rect 20404 21496 20410 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 21177 21539 21235 21545
rect 21177 21505 21189 21539
rect 21223 21536 21235 21539
rect 22646 21536 22652 21548
rect 21223 21508 22094 21536
rect 22607 21508 22652 21536
rect 21223 21505 21235 21508
rect 21177 21499 21235 21505
rect 15611 21372 17356 21400
rect 17431 21440 18828 21468
rect 15611 21369 15623 21372
rect 15565 21363 15623 21369
rect 3053 21335 3111 21341
rect 3053 21301 3065 21335
rect 3099 21332 3111 21335
rect 3234 21332 3240 21344
rect 3099 21304 3240 21332
rect 3099 21301 3111 21304
rect 3053 21295 3111 21301
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 9674 21332 9680 21344
rect 9635 21304 9680 21332
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 12253 21335 12311 21341
rect 12253 21301 12265 21335
rect 12299 21332 12311 21335
rect 12342 21332 12348 21344
rect 12299 21304 12348 21332
rect 12299 21301 12311 21304
rect 12253 21295 12311 21301
rect 12342 21292 12348 21304
rect 12400 21292 12406 21344
rect 13170 21332 13176 21344
rect 13131 21304 13176 21332
rect 13170 21292 13176 21304
rect 13228 21292 13234 21344
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 13357 21335 13415 21341
rect 13357 21332 13369 21335
rect 13320 21304 13369 21332
rect 13320 21292 13326 21304
rect 13357 21301 13369 21304
rect 13403 21301 13415 21335
rect 13357 21295 13415 21301
rect 14921 21335 14979 21341
rect 14921 21301 14933 21335
rect 14967 21332 14979 21335
rect 15838 21332 15844 21344
rect 14967 21304 15844 21332
rect 14967 21301 14979 21304
rect 14921 21295 14979 21301
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 17431 21332 17459 21440
rect 17681 21403 17739 21409
rect 17681 21369 17693 21403
rect 17727 21400 17739 21403
rect 17770 21400 17776 21412
rect 17727 21372 17776 21400
rect 17727 21369 17739 21372
rect 17681 21363 17739 21369
rect 17770 21360 17776 21372
rect 17828 21400 17834 21412
rect 20254 21400 20260 21412
rect 17828 21372 20260 21400
rect 17828 21360 17834 21372
rect 20254 21360 20260 21372
rect 20312 21400 20318 21412
rect 21910 21400 21916 21412
rect 20312 21372 21916 21400
rect 20312 21360 20318 21372
rect 21910 21360 21916 21372
rect 21968 21360 21974 21412
rect 17184 21304 17459 21332
rect 17497 21335 17555 21341
rect 17184 21292 17190 21304
rect 17497 21301 17509 21335
rect 17543 21332 17555 21335
rect 18230 21332 18236 21344
rect 17543 21304 18236 21332
rect 17543 21301 17555 21304
rect 17497 21295 17555 21301
rect 18230 21292 18236 21304
rect 18288 21332 18294 21344
rect 18782 21332 18788 21344
rect 18288 21304 18788 21332
rect 18288 21292 18294 21304
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 18877 21335 18935 21341
rect 18877 21301 18889 21335
rect 18923 21332 18935 21335
rect 19334 21332 19340 21344
rect 18923 21304 19340 21332
rect 18923 21301 18935 21304
rect 18877 21295 18935 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 22066 21332 22094 21508
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 23750 21536 23756 21548
rect 23711 21508 23756 21536
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 23934 21536 23940 21548
rect 23895 21508 23940 21536
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24044 21545 24072 21576
rect 27154 21564 27160 21576
rect 27212 21564 27218 21616
rect 35434 21604 35440 21616
rect 35395 21576 35440 21604
rect 35434 21564 35440 21576
rect 35492 21564 35498 21616
rect 24029 21539 24087 21545
rect 24029 21505 24041 21539
rect 24075 21505 24087 21539
rect 24029 21499 24087 21505
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 26694 21536 26700 21548
rect 24176 21508 26700 21536
rect 24176 21496 24182 21508
rect 26694 21496 26700 21508
rect 26752 21496 26758 21548
rect 27706 21536 27712 21548
rect 27667 21508 27712 21536
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 27982 21545 27988 21548
rect 27976 21536 27988 21545
rect 27943 21508 27988 21536
rect 27976 21499 27988 21508
rect 27982 21496 27988 21499
rect 28040 21496 28046 21548
rect 29546 21536 29552 21548
rect 29507 21508 29552 21536
rect 29546 21496 29552 21508
rect 29604 21496 29610 21548
rect 29733 21539 29791 21545
rect 29733 21505 29745 21539
rect 29779 21536 29791 21539
rect 30374 21536 30380 21548
rect 29779 21508 30380 21536
rect 29779 21505 29791 21508
rect 29733 21499 29791 21505
rect 30374 21496 30380 21508
rect 30432 21496 30438 21548
rect 32950 21536 32956 21548
rect 32911 21508 32956 21536
rect 32950 21496 32956 21508
rect 33008 21496 33014 21548
rect 33594 21536 33600 21548
rect 33555 21508 33600 21536
rect 33594 21496 33600 21508
rect 33652 21496 33658 21548
rect 22741 21471 22799 21477
rect 22741 21437 22753 21471
rect 22787 21468 22799 21471
rect 23566 21468 23572 21480
rect 22787 21440 23572 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 33045 21471 33103 21477
rect 33045 21437 33057 21471
rect 33091 21468 33103 21471
rect 33781 21471 33839 21477
rect 33781 21468 33793 21471
rect 33091 21440 33793 21468
rect 33091 21437 33103 21440
rect 33045 21431 33103 21437
rect 33781 21437 33793 21440
rect 33827 21437 33839 21471
rect 33781 21431 33839 21437
rect 23017 21403 23075 21409
rect 23017 21369 23029 21403
rect 23063 21400 23075 21403
rect 23658 21400 23664 21412
rect 23063 21372 23664 21400
rect 23063 21369 23075 21372
rect 23017 21363 23075 21369
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 27430 21332 27436 21344
rect 22066 21304 27436 21332
rect 27430 21292 27436 21304
rect 27488 21292 27494 21344
rect 28442 21292 28448 21344
rect 28500 21332 28506 21344
rect 29089 21335 29147 21341
rect 29089 21332 29101 21335
rect 28500 21304 29101 21332
rect 28500 21292 28506 21304
rect 29089 21301 29101 21304
rect 29135 21301 29147 21335
rect 29089 21295 29147 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 8389 21131 8447 21137
rect 8389 21097 8401 21131
rect 8435 21128 8447 21131
rect 9122 21128 9128 21140
rect 8435 21100 9128 21128
rect 8435 21097 8447 21100
rect 8389 21091 8447 21097
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13541 21131 13599 21137
rect 13541 21128 13553 21131
rect 13228 21100 13553 21128
rect 13228 21088 13234 21100
rect 13541 21097 13553 21100
rect 13587 21097 13599 21131
rect 13541 21091 13599 21097
rect 17129 21131 17187 21137
rect 17129 21097 17141 21131
rect 17175 21128 17187 21131
rect 17402 21128 17408 21140
rect 17175 21100 17408 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 17402 21088 17408 21100
rect 17460 21088 17466 21140
rect 24854 21128 24860 21140
rect 24596 21100 24860 21128
rect 14829 21063 14887 21069
rect 14829 21029 14841 21063
rect 14875 21060 14887 21063
rect 20070 21060 20076 21072
rect 14875 21032 20076 21060
rect 14875 21029 14887 21032
rect 14829 21023 14887 21029
rect 20070 21020 20076 21032
rect 20128 21020 20134 21072
rect 22094 21020 22100 21072
rect 22152 21020 22158 21072
rect 1578 20992 1584 21004
rect 1539 20964 1584 20992
rect 1578 20952 1584 20964
rect 1636 20952 1642 21004
rect 3234 20992 3240 21004
rect 3195 20964 3240 20992
rect 3234 20952 3240 20964
rect 3292 20952 3298 21004
rect 8573 20995 8631 21001
rect 8573 20961 8585 20995
rect 8619 20961 8631 20995
rect 8573 20955 8631 20961
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 8294 20924 8300 20936
rect 8255 20896 8300 20924
rect 3421 20887 3479 20893
rect 3050 20816 3056 20868
rect 3108 20856 3114 20868
rect 3436 20856 3464 20887
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 3108 20828 3464 20856
rect 8588 20856 8616 20955
rect 8662 20952 8668 21004
rect 8720 20992 8726 21004
rect 9493 20995 9551 21001
rect 9493 20992 9505 20995
rect 8720 20964 9505 20992
rect 8720 20952 8726 20964
rect 9493 20961 9505 20964
rect 9539 20961 9551 20995
rect 9493 20955 9551 20961
rect 13446 20952 13452 21004
rect 13504 20992 13510 21004
rect 14553 20995 14611 21001
rect 14553 20992 14565 20995
rect 13504 20964 14565 20992
rect 13504 20952 13510 20964
rect 14553 20961 14565 20964
rect 14599 20961 14611 20995
rect 14553 20955 14611 20961
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 18782 20992 18788 21004
rect 14700 20964 18788 20992
rect 14700 20952 14706 20964
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 22112 20992 22140 21020
rect 24596 21001 24624 21100
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 27982 21128 27988 21140
rect 27943 21100 27988 21128
rect 27982 21088 27988 21100
rect 28040 21088 28046 21140
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 22112 20964 22569 20992
rect 22557 20961 22569 20964
rect 22603 20992 22615 20995
rect 24581 20995 24639 21001
rect 24581 20992 24593 20995
rect 22603 20964 24593 20992
rect 22603 20961 22615 20964
rect 22557 20955 22615 20961
rect 24581 20961 24593 20964
rect 24627 20961 24639 20995
rect 24581 20955 24639 20961
rect 26234 20952 26240 21004
rect 26292 20992 26298 21004
rect 26421 20995 26479 21001
rect 26421 20992 26433 20995
rect 26292 20964 26433 20992
rect 26292 20952 26298 20964
rect 26421 20961 26433 20964
rect 26467 20961 26479 20995
rect 26694 20992 26700 21004
rect 26655 20964 26700 20992
rect 26421 20955 26479 20961
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 8846 20884 8852 20936
rect 8904 20924 8910 20936
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 8904 20896 9321 20924
rect 8904 20884 8910 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20924 10379 20927
rect 12158 20924 12164 20936
rect 10367 20896 12164 20924
rect 10367 20893 10379 20896
rect 10321 20887 10379 20893
rect 10704 20868 10732 20896
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 14366 20924 14372 20936
rect 14327 20896 14372 20924
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 17218 20924 17224 20936
rect 14516 20896 14561 20924
rect 17179 20896 17224 20924
rect 14516 20884 14522 20896
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 17586 20884 17592 20936
rect 17644 20924 17650 20936
rect 17865 20927 17923 20933
rect 17865 20924 17877 20927
rect 17644 20896 17877 20924
rect 17644 20884 17650 20896
rect 17865 20893 17877 20896
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20924 18107 20927
rect 18506 20924 18512 20936
rect 18095 20896 18512 20924
rect 18095 20893 18107 20896
rect 18049 20887 18107 20893
rect 9582 20856 9588 20868
rect 8588 20828 9588 20856
rect 3108 20816 3114 20828
rect 9582 20816 9588 20828
rect 9640 20816 9646 20868
rect 9674 20816 9680 20868
rect 9732 20856 9738 20868
rect 10566 20859 10624 20865
rect 10566 20856 10578 20859
rect 9732 20828 10578 20856
rect 9732 20816 9738 20828
rect 10566 20825 10578 20828
rect 10612 20825 10624 20859
rect 10566 20819 10624 20825
rect 10686 20816 10692 20868
rect 10744 20816 10750 20868
rect 12434 20865 12440 20868
rect 12428 20819 12440 20865
rect 12492 20856 12498 20868
rect 17880 20856 17908 20887
rect 18506 20884 18512 20896
rect 18564 20884 18570 20936
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20924 19671 20927
rect 19978 20924 19984 20936
rect 19659 20896 19984 20924
rect 19659 20893 19671 20896
rect 19613 20887 19671 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 20806 20924 20812 20936
rect 20767 20896 20812 20924
rect 20806 20884 20812 20896
rect 20864 20924 20870 20936
rect 22094 20924 22100 20936
rect 20864 20896 22100 20924
rect 20864 20884 20870 20896
rect 22094 20884 22100 20896
rect 22152 20884 22158 20936
rect 23382 20884 23388 20936
rect 23440 20924 23446 20936
rect 24837 20927 24895 20933
rect 24837 20924 24849 20927
rect 23440 20896 24849 20924
rect 23440 20884 23446 20896
rect 24837 20893 24849 20896
rect 24883 20893 24895 20927
rect 27706 20924 27712 20936
rect 27667 20896 27712 20924
rect 24837 20887 24895 20893
rect 27706 20884 27712 20896
rect 27764 20884 27770 20936
rect 28442 20924 28448 20936
rect 27816 20896 28448 20924
rect 18693 20859 18751 20865
rect 18693 20856 18705 20859
rect 12492 20828 12528 20856
rect 17880 20828 18705 20856
rect 12434 20816 12440 20819
rect 12492 20816 12498 20828
rect 18693 20825 18705 20828
rect 18739 20825 18751 20859
rect 18693 20819 18751 20825
rect 19794 20816 19800 20868
rect 19852 20856 19858 20868
rect 26602 20856 26608 20868
rect 19852 20828 26608 20856
rect 19852 20816 19858 20828
rect 26602 20816 26608 20828
rect 26660 20856 26666 20868
rect 27816 20856 27844 20896
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28626 20924 28632 20936
rect 28587 20896 28632 20924
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 26660 20828 27844 20856
rect 26660 20816 26666 20828
rect 27890 20816 27896 20868
rect 27948 20856 27954 20868
rect 27985 20859 28043 20865
rect 27985 20856 27997 20859
rect 27948 20828 27997 20856
rect 27948 20816 27954 20828
rect 27985 20825 27997 20828
rect 28031 20856 28043 20859
rect 28166 20856 28172 20868
rect 28031 20828 28172 20856
rect 28031 20825 28043 20828
rect 27985 20819 28043 20825
rect 28166 20816 28172 20828
rect 28224 20816 28230 20868
rect 8570 20788 8576 20800
rect 8531 20760 8576 20788
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 11701 20791 11759 20797
rect 11701 20757 11713 20791
rect 11747 20788 11759 20791
rect 12986 20788 12992 20800
rect 11747 20760 12992 20788
rect 11747 20757 11759 20760
rect 11701 20751 11759 20757
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 16758 20748 16764 20800
rect 16816 20788 16822 20800
rect 17034 20788 17040 20800
rect 16816 20760 17040 20788
rect 16816 20748 16822 20760
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17954 20788 17960 20800
rect 17915 20760 17960 20788
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 18877 20791 18935 20797
rect 18877 20757 18889 20791
rect 18923 20788 18935 20791
rect 18966 20788 18972 20800
rect 18923 20760 18972 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 18966 20748 18972 20760
rect 19024 20748 19030 20800
rect 19426 20788 19432 20800
rect 19387 20760 19432 20788
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 25961 20791 26019 20797
rect 25961 20757 25973 20791
rect 26007 20788 26019 20791
rect 26326 20788 26332 20800
rect 26007 20760 26332 20788
rect 26007 20757 26019 20760
rect 25961 20751 26019 20757
rect 26326 20748 26332 20760
rect 26384 20748 26390 20800
rect 27801 20791 27859 20797
rect 27801 20757 27813 20791
rect 27847 20788 27859 20791
rect 28445 20791 28503 20797
rect 28445 20788 28457 20791
rect 27847 20760 28457 20788
rect 27847 20757 27859 20760
rect 27801 20751 27859 20757
rect 28445 20757 28457 20760
rect 28491 20757 28503 20791
rect 28445 20751 28503 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 8957 20587 9015 20593
rect 8957 20584 8969 20587
rect 8904 20556 8969 20584
rect 8904 20544 8910 20556
rect 8957 20553 8969 20556
rect 9003 20553 9015 20587
rect 8957 20547 9015 20553
rect 9677 20587 9735 20593
rect 9677 20553 9689 20587
rect 9723 20584 9735 20587
rect 12434 20584 12440 20596
rect 9723 20556 12440 20584
rect 9723 20553 9735 20556
rect 9677 20547 9735 20553
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 13633 20587 13691 20593
rect 13633 20553 13645 20587
rect 13679 20584 13691 20587
rect 16758 20584 16764 20596
rect 13679 20556 16764 20584
rect 13679 20553 13691 20556
rect 13633 20547 13691 20553
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 16942 20584 16948 20596
rect 16903 20556 16948 20584
rect 16942 20544 16948 20556
rect 17000 20584 17006 20596
rect 17402 20584 17408 20596
rect 17000 20556 17408 20584
rect 17000 20544 17006 20556
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 20073 20587 20131 20593
rect 20073 20553 20085 20587
rect 20119 20584 20131 20587
rect 20806 20584 20812 20596
rect 20119 20556 20812 20584
rect 20119 20553 20131 20556
rect 20073 20547 20131 20553
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 27325 20587 27383 20593
rect 27325 20584 27337 20587
rect 26436 20556 27337 20584
rect 1946 20516 1952 20528
rect 1907 20488 1952 20516
rect 1946 20476 1952 20488
rect 2004 20476 2010 20528
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 8757 20519 8815 20525
rect 8757 20516 8769 20519
rect 8352 20488 8769 20516
rect 8352 20476 8358 20488
rect 8757 20485 8769 20488
rect 8803 20516 8815 20519
rect 13170 20516 13176 20528
rect 8803 20488 12434 20516
rect 8803 20485 8815 20488
rect 8757 20479 8815 20485
rect 8570 20408 8576 20460
rect 8628 20448 8634 20460
rect 9585 20451 9643 20457
rect 9585 20448 9597 20451
rect 8628 20420 9597 20448
rect 8628 20408 8634 20420
rect 9585 20417 9597 20420
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20417 9827 20451
rect 9769 20411 9827 20417
rect 2682 20340 2688 20392
rect 2740 20380 2746 20392
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 2740 20352 3617 20380
rect 2740 20340 2746 20352
rect 3605 20349 3617 20352
rect 3651 20349 3663 20383
rect 3786 20380 3792 20392
rect 3747 20352 3792 20380
rect 3605 20343 3663 20349
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 9784 20380 9812 20411
rect 9140 20352 9812 20380
rect 9140 20324 9168 20352
rect 9122 20312 9128 20324
rect 9035 20284 9128 20312
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 12406 20312 12434 20488
rect 12820 20488 13176 20516
rect 12820 20457 12848 20488
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 17954 20476 17960 20528
rect 18012 20516 18018 20528
rect 19153 20519 19211 20525
rect 19153 20516 19165 20519
rect 18012 20488 19165 20516
rect 18012 20476 18018 20488
rect 19153 20485 19165 20488
rect 19199 20485 19211 20519
rect 19153 20479 19211 20485
rect 19245 20519 19303 20525
rect 19245 20485 19257 20519
rect 19291 20516 19303 20519
rect 19426 20516 19432 20528
rect 19291 20488 19432 20516
rect 19291 20485 19303 20488
rect 19245 20479 19303 20485
rect 19426 20476 19432 20488
rect 19484 20476 19490 20528
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 13262 20448 13268 20460
rect 13223 20420 13268 20448
rect 12805 20411 12863 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13906 20408 13912 20460
rect 13964 20448 13970 20460
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 13964 20420 14933 20448
rect 13964 20408 13970 20420
rect 14921 20417 14933 20420
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20448 16911 20451
rect 17586 20448 17592 20460
rect 16899 20420 17592 20448
rect 16899 20417 16911 20420
rect 16853 20411 16911 20417
rect 14936 20380 14964 20411
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20417 17739 20451
rect 18966 20448 18972 20460
rect 18927 20420 18972 20448
rect 17681 20411 17739 20417
rect 17696 20380 17724 20411
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 19334 20448 19340 20460
rect 19295 20420 19340 20448
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 21174 20448 21180 20460
rect 21232 20457 21238 20460
rect 21144 20420 21180 20448
rect 21174 20408 21180 20420
rect 21232 20411 21244 20457
rect 21453 20451 21511 20457
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 22002 20448 22008 20460
rect 21499 20420 22008 20448
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 21232 20408 21238 20411
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 22278 20448 22284 20460
rect 22239 20420 22284 20448
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 26234 20408 26240 20460
rect 26292 20448 26298 20460
rect 26436 20457 26464 20556
rect 27325 20553 27337 20556
rect 27371 20584 27383 20587
rect 30558 20584 30564 20596
rect 27371 20556 28304 20584
rect 30519 20556 30564 20584
rect 27371 20553 27383 20556
rect 27325 20547 27383 20553
rect 26694 20476 26700 20528
rect 26752 20516 26758 20528
rect 27525 20519 27583 20525
rect 27525 20516 27537 20519
rect 26752 20488 27537 20516
rect 26752 20476 26758 20488
rect 27525 20485 27537 20488
rect 27571 20516 27583 20519
rect 27985 20519 28043 20525
rect 27985 20516 27997 20519
rect 27571 20488 27997 20516
rect 27571 20485 27583 20488
rect 27525 20479 27583 20485
rect 27985 20485 27997 20488
rect 28031 20485 28043 20519
rect 27985 20479 28043 20485
rect 26329 20451 26387 20457
rect 26329 20448 26341 20451
rect 26292 20420 26341 20448
rect 26292 20408 26298 20420
rect 26329 20417 26341 20420
rect 26375 20417 26387 20451
rect 26329 20411 26387 20417
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20448 26479 20451
rect 26510 20448 26516 20460
rect 26467 20420 26516 20448
rect 26467 20417 26479 20420
rect 26421 20411 26479 20417
rect 26510 20408 26516 20420
rect 26568 20408 26574 20460
rect 26605 20451 26663 20457
rect 26605 20417 26617 20451
rect 26651 20448 26663 20451
rect 28074 20448 28080 20460
rect 26651 20420 28080 20448
rect 26651 20417 26663 20420
rect 26605 20411 26663 20417
rect 28074 20408 28080 20420
rect 28132 20408 28138 20460
rect 28276 20457 28304 20556
rect 30558 20544 30564 20556
rect 30616 20584 30622 20596
rect 30926 20584 30932 20596
rect 30616 20556 30932 20584
rect 30616 20544 30622 20556
rect 30926 20544 30932 20556
rect 30984 20544 30990 20596
rect 28169 20451 28227 20457
rect 28169 20417 28181 20451
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 28261 20451 28319 20457
rect 28261 20417 28273 20451
rect 28307 20417 28319 20451
rect 28261 20411 28319 20417
rect 19978 20380 19984 20392
rect 14936 20352 19984 20380
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 22373 20383 22431 20389
rect 22373 20349 22385 20383
rect 22419 20380 22431 20383
rect 24026 20380 24032 20392
rect 22419 20352 24032 20380
rect 22419 20349 22431 20352
rect 22373 20343 22431 20349
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20349 26019 20383
rect 27890 20380 27896 20392
rect 25961 20343 26019 20349
rect 27356 20352 27896 20380
rect 12621 20315 12679 20321
rect 12621 20312 12633 20315
rect 12406 20284 12633 20312
rect 12621 20281 12633 20284
rect 12667 20312 12679 20315
rect 17954 20312 17960 20324
rect 12667 20284 17960 20312
rect 12667 20281 12679 20284
rect 12621 20275 12679 20281
rect 17954 20272 17960 20284
rect 18012 20272 18018 20324
rect 19521 20315 19579 20321
rect 19521 20281 19533 20315
rect 19567 20312 19579 20315
rect 22649 20315 22707 20321
rect 19567 20284 20576 20312
rect 19567 20281 19579 20284
rect 19521 20275 19579 20281
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 8720 20216 8953 20244
rect 8720 20204 8726 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 8941 20207 8999 20213
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13449 20247 13507 20253
rect 13449 20244 13461 20247
rect 13136 20216 13461 20244
rect 13136 20204 13142 20216
rect 13449 20213 13461 20216
rect 13495 20244 13507 20247
rect 14642 20244 14648 20256
rect 13495 20216 14648 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 14642 20204 14648 20216
rect 14700 20204 14706 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 15013 20247 15071 20253
rect 15013 20244 15025 20247
rect 14884 20216 15025 20244
rect 14884 20204 14890 20216
rect 15013 20213 15025 20216
rect 15059 20244 15071 20247
rect 17126 20244 17132 20256
rect 15059 20216 17132 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17310 20204 17316 20256
rect 17368 20244 17374 20256
rect 17589 20247 17647 20253
rect 17589 20244 17601 20247
rect 17368 20216 17601 20244
rect 17368 20204 17374 20216
rect 17589 20213 17601 20216
rect 17635 20213 17647 20247
rect 20548 20244 20576 20284
rect 22649 20281 22661 20315
rect 22695 20312 22707 20315
rect 23198 20312 23204 20324
rect 22695 20284 23204 20312
rect 22695 20281 22707 20284
rect 22649 20275 22707 20281
rect 23198 20272 23204 20284
rect 23256 20272 23262 20324
rect 25976 20312 26004 20343
rect 27356 20312 27384 20352
rect 27890 20340 27896 20352
rect 27948 20380 27954 20392
rect 28184 20380 28212 20411
rect 30466 20408 30472 20460
rect 30524 20457 30530 20460
rect 30524 20451 30560 20457
rect 30548 20417 30560 20451
rect 30524 20411 30560 20417
rect 30524 20408 30530 20411
rect 31110 20408 31116 20460
rect 31168 20448 31174 20460
rect 31481 20451 31539 20457
rect 31481 20448 31493 20451
rect 31168 20420 31493 20448
rect 31168 20408 31174 20420
rect 31481 20417 31493 20420
rect 31527 20417 31539 20451
rect 31481 20411 31539 20417
rect 27948 20352 28212 20380
rect 31021 20383 31079 20389
rect 27948 20340 27954 20352
rect 31021 20349 31033 20383
rect 31067 20380 31079 20383
rect 31662 20380 31668 20392
rect 31067 20352 31668 20380
rect 31067 20349 31079 20352
rect 31021 20343 31079 20349
rect 31662 20340 31668 20352
rect 31720 20340 31726 20392
rect 25976 20284 27384 20312
rect 20714 20244 20720 20256
rect 20548 20216 20720 20244
rect 17589 20207 17647 20213
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 26970 20204 26976 20256
rect 27028 20244 27034 20256
rect 27356 20253 27384 20284
rect 30834 20272 30840 20324
rect 30892 20312 30898 20324
rect 31570 20312 31576 20324
rect 30892 20284 31576 20312
rect 30892 20272 30898 20284
rect 31570 20272 31576 20284
rect 31628 20272 31634 20324
rect 27157 20247 27215 20253
rect 27157 20244 27169 20247
rect 27028 20216 27169 20244
rect 27028 20204 27034 20216
rect 27157 20213 27169 20216
rect 27203 20213 27215 20247
rect 27157 20207 27215 20213
rect 27341 20247 27399 20253
rect 27341 20213 27353 20247
rect 27387 20213 27399 20247
rect 27982 20244 27988 20256
rect 27943 20216 27988 20244
rect 27341 20207 27399 20213
rect 27982 20204 27988 20216
rect 28040 20204 28046 20256
rect 29914 20204 29920 20256
rect 29972 20244 29978 20256
rect 30377 20247 30435 20253
rect 30377 20244 30389 20247
rect 29972 20216 30389 20244
rect 29972 20204 29978 20216
rect 30377 20213 30389 20216
rect 30423 20213 30435 20247
rect 30377 20207 30435 20213
rect 30558 20204 30564 20256
rect 30616 20244 30622 20256
rect 30742 20244 30748 20256
rect 30616 20216 30748 20244
rect 30616 20204 30622 20216
rect 30742 20204 30748 20216
rect 30800 20244 30806 20256
rect 30929 20247 30987 20253
rect 30929 20244 30941 20247
rect 30800 20216 30941 20244
rect 30800 20204 30806 20216
rect 30929 20213 30941 20216
rect 30975 20213 30987 20247
rect 30929 20207 30987 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2682 20040 2688 20052
rect 2643 20012 2688 20040
rect 2682 20000 2688 20012
rect 2740 20000 2746 20052
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 3786 20040 3792 20052
rect 3467 20012 3792 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 16298 20040 16304 20052
rect 14568 20012 16304 20040
rect 2133 19975 2191 19981
rect 2133 19941 2145 19975
rect 2179 19972 2191 19975
rect 3050 19972 3056 19984
rect 2179 19944 3056 19972
rect 2179 19941 2191 19944
rect 2133 19935 2191 19941
rect 3050 19932 3056 19944
rect 3108 19932 3114 19984
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19805 2835 19839
rect 2777 19799 2835 19805
rect 2792 19768 2820 19799
rect 4062 19796 4068 19848
rect 4120 19836 4126 19848
rect 5626 19836 5632 19848
rect 4120 19808 5632 19836
rect 4120 19796 4126 19808
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 11974 19796 11980 19848
rect 12032 19836 12038 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 12032 19808 14289 19836
rect 12032 19796 12038 19808
rect 14277 19805 14289 19808
rect 14323 19836 14335 19839
rect 14458 19836 14464 19848
rect 14323 19808 14464 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 4706 19768 4712 19780
rect 2792 19740 4712 19768
rect 4706 19728 4712 19740
rect 4764 19768 4770 19780
rect 14568 19768 14596 20012
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 18196 20012 18337 20040
rect 18196 20000 18202 20012
rect 18325 20009 18337 20012
rect 18371 20009 18383 20043
rect 18325 20003 18383 20009
rect 20625 20043 20683 20049
rect 20625 20009 20637 20043
rect 20671 20009 20683 20043
rect 20625 20003 20683 20009
rect 16850 19932 16856 19984
rect 16908 19972 16914 19984
rect 20640 19972 20668 20003
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 21232 20012 21281 20040
rect 21232 20000 21238 20012
rect 21269 20009 21281 20012
rect 21315 20009 21327 20043
rect 21269 20003 21327 20009
rect 26421 20043 26479 20049
rect 26421 20009 26433 20043
rect 26467 20040 26479 20043
rect 26510 20040 26516 20052
rect 26467 20012 26516 20040
rect 26467 20009 26479 20012
rect 26421 20003 26479 20009
rect 26510 20000 26516 20012
rect 26568 20000 26574 20052
rect 27157 20043 27215 20049
rect 27157 20009 27169 20043
rect 27203 20040 27215 20043
rect 27982 20040 27988 20052
rect 27203 20012 27988 20040
rect 27203 20009 27215 20012
rect 27157 20003 27215 20009
rect 27982 20000 27988 20012
rect 28040 20000 28046 20052
rect 31110 20040 31116 20052
rect 31071 20012 31116 20040
rect 31110 20000 31116 20012
rect 31168 20000 31174 20052
rect 31662 20040 31668 20052
rect 31623 20012 31668 20040
rect 31662 20000 31668 20012
rect 31720 20000 31726 20052
rect 27341 19975 27399 19981
rect 16908 19944 17264 19972
rect 20640 19944 22094 19972
rect 16908 19932 16914 19944
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 16390 19904 16396 19916
rect 15335 19876 16396 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 17120 19904 17126 19916
rect 17081 19876 17126 19904
rect 17120 19864 17126 19876
rect 17178 19864 17184 19916
rect 17236 19913 17264 19944
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 15194 19836 15200 19848
rect 15155 19808 15200 19836
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 17037 19839 17095 19845
rect 15580 19826 16810 19836
rect 16841 19829 16899 19835
rect 16841 19826 16853 19829
rect 15580 19808 16853 19826
rect 4764 19740 14596 19768
rect 4764 19728 4770 19740
rect 10226 19660 10232 19712
rect 10284 19700 10290 19712
rect 14458 19700 14464 19712
rect 10284 19672 14464 19700
rect 10284 19660 10290 19672
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 15580 19709 15608 19808
rect 16782 19798 16853 19808
rect 16841 19795 16853 19798
rect 16887 19795 16899 19829
rect 17037 19805 17049 19839
rect 17083 19838 17095 19839
rect 17083 19814 17096 19838
rect 17402 19836 17408 19848
rect 17083 19805 17166 19814
rect 17363 19808 17408 19836
rect 17037 19799 17166 19805
rect 16841 19789 16899 19795
rect 17068 19786 17166 19799
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 20257 19839 20315 19845
rect 18748 19808 18793 19836
rect 18748 19796 18754 19808
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20714 19836 20720 19848
rect 20303 19808 20720 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 20714 19796 20720 19808
rect 20772 19836 20778 19848
rect 20990 19836 20996 19848
rect 20772 19808 20996 19836
rect 20772 19796 20778 19808
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21450 19836 21456 19848
rect 21411 19808 21456 19836
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 22066 19836 22094 19944
rect 27341 19941 27353 19975
rect 27387 19972 27399 19975
rect 27706 19972 27712 19984
rect 27387 19944 27712 19972
rect 27387 19941 27399 19944
rect 27341 19935 27399 19941
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 27890 19972 27896 19984
rect 27851 19944 27896 19972
rect 27890 19932 27896 19944
rect 27948 19932 27954 19984
rect 26602 19904 26608 19916
rect 26068 19876 26608 19904
rect 23658 19836 23664 19848
rect 22066 19808 23664 19836
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 24026 19836 24032 19848
rect 23987 19808 24032 19836
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 26068 19845 26096 19876
rect 26602 19864 26608 19876
rect 26660 19904 26666 19916
rect 26660 19876 28028 19904
rect 26660 19864 26666 19876
rect 26053 19839 26111 19845
rect 26053 19805 26065 19839
rect 26099 19805 26111 19839
rect 26053 19799 26111 19805
rect 26237 19839 26295 19845
rect 26237 19805 26249 19839
rect 26283 19836 26295 19839
rect 26326 19836 26332 19848
rect 26283 19808 26332 19836
rect 26283 19805 26295 19808
rect 26237 19799 26295 19805
rect 26326 19796 26332 19808
rect 26384 19796 26390 19848
rect 26970 19836 26976 19848
rect 26931 19808 26976 19836
rect 26970 19796 26976 19808
rect 27028 19796 27034 19848
rect 27154 19836 27160 19848
rect 27115 19808 27160 19836
rect 27154 19796 27160 19808
rect 27212 19836 27218 19848
rect 27522 19836 27528 19848
rect 27212 19808 27528 19836
rect 27212 19796 27218 19808
rect 27522 19796 27528 19808
rect 27580 19796 27586 19848
rect 27614 19796 27620 19848
rect 27672 19836 27678 19848
rect 28000 19845 28028 19876
rect 30098 19864 30104 19916
rect 30156 19904 30162 19916
rect 30653 19907 30711 19913
rect 30653 19904 30665 19907
rect 30156 19876 30665 19904
rect 30156 19864 30162 19876
rect 30653 19873 30665 19876
rect 30699 19873 30711 19907
rect 31846 19904 31852 19916
rect 31807 19876 31852 19904
rect 30653 19867 30711 19873
rect 31846 19864 31852 19876
rect 31904 19864 31910 19916
rect 27801 19839 27859 19845
rect 27801 19836 27813 19839
rect 27672 19808 27813 19836
rect 27672 19796 27678 19808
rect 27801 19805 27813 19808
rect 27847 19805 27859 19839
rect 27801 19799 27859 19805
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19805 28043 19839
rect 27985 19799 28043 19805
rect 29086 19796 29092 19848
rect 29144 19836 29150 19848
rect 29546 19836 29552 19848
rect 29144 19808 29552 19836
rect 29144 19796 29150 19808
rect 29546 19796 29552 19808
rect 29604 19836 29610 19848
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29604 19808 29745 19836
rect 29604 19796 29610 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29914 19836 29920 19848
rect 29875 19808 29920 19836
rect 29733 19799 29791 19805
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 30745 19839 30803 19845
rect 30745 19805 30757 19839
rect 30791 19805 30803 19839
rect 30745 19799 30803 19805
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 16117 19771 16175 19777
rect 16117 19768 16129 19771
rect 15896 19740 16129 19768
rect 15896 19728 15902 19740
rect 16117 19737 16129 19740
rect 16163 19737 16175 19771
rect 17138 19768 17166 19786
rect 18322 19768 18328 19780
rect 17138 19740 18328 19768
rect 16117 19731 16175 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 18874 19768 18880 19780
rect 18835 19740 18880 19768
rect 18874 19728 18880 19740
rect 18932 19768 18938 19780
rect 19426 19768 19432 19780
rect 18932 19740 19432 19768
rect 18932 19728 18938 19740
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 22186 19768 22192 19780
rect 19536 19740 22192 19768
rect 15565 19703 15623 19709
rect 15565 19669 15577 19703
rect 15611 19669 15623 19703
rect 15565 19663 15623 19669
rect 15930 19660 15936 19712
rect 15988 19700 15994 19712
rect 16209 19703 16267 19709
rect 16209 19700 16221 19703
rect 15988 19672 16221 19700
rect 15988 19660 15994 19672
rect 16209 19669 16221 19672
rect 16255 19700 16267 19703
rect 16666 19700 16672 19712
rect 16255 19672 16672 19700
rect 16255 19669 16267 19672
rect 16209 19663 16267 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 17126 19660 17132 19712
rect 17184 19700 17190 19712
rect 17589 19703 17647 19709
rect 17589 19700 17601 19703
rect 17184 19672 17601 19700
rect 17184 19660 17190 19672
rect 17589 19669 17601 19672
rect 17635 19669 17647 19703
rect 17589 19663 17647 19669
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18012 19672 18521 19700
rect 18012 19660 18018 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 18782 19700 18788 19712
rect 18647 19672 18788 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 18782 19660 18788 19672
rect 18840 19700 18846 19712
rect 19536 19700 19564 19740
rect 22186 19728 22192 19740
rect 22244 19768 22250 19780
rect 22646 19768 22652 19780
rect 22244 19740 22652 19768
rect 22244 19728 22250 19740
rect 22646 19728 22652 19740
rect 22704 19728 22710 19780
rect 23753 19771 23811 19777
rect 23753 19737 23765 19771
rect 23799 19737 23811 19771
rect 23753 19731 23811 19737
rect 23845 19771 23903 19777
rect 23845 19737 23857 19771
rect 23891 19768 23903 19771
rect 24118 19768 24124 19780
rect 23891 19740 24124 19768
rect 23891 19737 23903 19740
rect 23845 19731 23903 19737
rect 18840 19672 19564 19700
rect 18840 19660 18846 19672
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20625 19703 20683 19709
rect 20625 19700 20637 19703
rect 20036 19672 20637 19700
rect 20036 19660 20042 19672
rect 20625 19669 20637 19672
rect 20671 19669 20683 19703
rect 20625 19663 20683 19669
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 20809 19703 20867 19709
rect 20809 19700 20821 19703
rect 20772 19672 20821 19700
rect 20772 19660 20778 19672
rect 20809 19669 20821 19672
rect 20855 19669 20867 19703
rect 20809 19663 20867 19669
rect 23477 19703 23535 19709
rect 23477 19669 23489 19703
rect 23523 19700 23535 19703
rect 23566 19700 23572 19712
rect 23523 19672 23572 19700
rect 23523 19669 23535 19672
rect 23477 19663 23535 19669
rect 23566 19660 23572 19672
rect 23624 19660 23630 19712
rect 23768 19700 23796 19731
rect 24118 19728 24124 19740
rect 24176 19728 24182 19780
rect 26344 19768 26372 19796
rect 30650 19768 30656 19780
rect 26344 19740 30656 19768
rect 30650 19728 30656 19740
rect 30708 19768 30714 19780
rect 30760 19768 30788 19799
rect 31570 19796 31576 19848
rect 31628 19836 31634 19848
rect 31941 19839 31999 19845
rect 31941 19836 31953 19839
rect 31628 19808 31953 19836
rect 31628 19796 31634 19808
rect 31941 19805 31953 19808
rect 31987 19805 31999 19839
rect 31941 19799 31999 19805
rect 37366 19796 37372 19848
rect 37424 19836 37430 19848
rect 37461 19839 37519 19845
rect 37461 19836 37473 19839
rect 37424 19808 37473 19836
rect 37424 19796 37430 19808
rect 37461 19805 37473 19808
rect 37507 19805 37519 19839
rect 37461 19799 37519 19805
rect 30708 19740 30788 19768
rect 30708 19728 30714 19740
rect 24486 19700 24492 19712
rect 23768 19672 24492 19700
rect 24486 19660 24492 19672
rect 24544 19660 24550 19712
rect 29822 19700 29828 19712
rect 29783 19672 29828 19700
rect 29822 19660 29828 19672
rect 29880 19660 29886 19712
rect 37553 19703 37611 19709
rect 37553 19669 37565 19703
rect 37599 19700 37611 19703
rect 38102 19700 38108 19712
rect 37599 19672 38108 19700
rect 37599 19669 37611 19672
rect 37553 19663 37611 19669
rect 38102 19660 38108 19672
rect 38160 19660 38166 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 9876 19468 12434 19496
rect 2777 19431 2835 19437
rect 2777 19397 2789 19431
rect 2823 19428 2835 19431
rect 3050 19428 3056 19440
rect 2823 19400 3056 19428
rect 2823 19397 2835 19400
rect 2777 19391 2835 19397
rect 3050 19388 3056 19400
rect 3108 19428 3114 19440
rect 3878 19428 3884 19440
rect 3108 19400 3884 19428
rect 3108 19388 3114 19400
rect 3878 19388 3884 19400
rect 3936 19388 3942 19440
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 3970 19360 3976 19372
rect 2547 19332 3976 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 3970 19320 3976 19332
rect 4028 19360 4034 19372
rect 9876 19369 9904 19468
rect 10505 19431 10563 19437
rect 10505 19397 10517 19431
rect 10551 19428 10563 19431
rect 11054 19428 11060 19440
rect 10551 19400 11060 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 12406 19428 12434 19468
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 13541 19499 13599 19505
rect 13541 19496 13553 19499
rect 13504 19468 13553 19496
rect 13504 19456 13510 19468
rect 13541 19465 13553 19468
rect 13587 19465 13599 19499
rect 17126 19496 17132 19508
rect 17087 19468 17132 19496
rect 13541 19459 13599 19465
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 18322 19496 18328 19508
rect 18283 19468 18328 19496
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 20073 19499 20131 19505
rect 20073 19465 20085 19499
rect 20119 19496 20131 19499
rect 21450 19496 21456 19508
rect 20119 19468 21456 19496
rect 20119 19465 20131 19468
rect 20073 19459 20131 19465
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 30098 19496 30104 19508
rect 27264 19468 30104 19496
rect 15286 19428 15292 19440
rect 12406 19400 15292 19428
rect 15286 19388 15292 19400
rect 15344 19388 15350 19440
rect 17218 19428 17224 19440
rect 16040 19400 17224 19428
rect 16040 19372 16068 19400
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 17678 19428 17684 19440
rect 17639 19400 17684 19428
rect 17678 19388 17684 19400
rect 17736 19388 17742 19440
rect 19334 19388 19340 19440
rect 19392 19428 19398 19440
rect 19705 19431 19763 19437
rect 19705 19428 19717 19431
rect 19392 19400 19717 19428
rect 19392 19388 19398 19400
rect 19705 19397 19717 19400
rect 19751 19397 19763 19431
rect 19705 19391 19763 19397
rect 19921 19431 19979 19437
rect 19921 19397 19933 19431
rect 19967 19428 19979 19431
rect 20162 19428 20168 19440
rect 19967 19400 20168 19428
rect 19967 19397 19979 19400
rect 19921 19391 19979 19397
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 20806 19388 20812 19440
rect 20864 19428 20870 19440
rect 20864 19400 21036 19428
rect 20864 19388 20870 19400
rect 4065 19363 4123 19369
rect 4065 19360 4077 19363
rect 4028 19332 4077 19360
rect 4028 19320 4034 19332
rect 4065 19329 4077 19332
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19329 9919 19363
rect 9861 19323 9919 19329
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 10137 19363 10195 19369
rect 10137 19329 10149 19363
rect 10183 19329 10195 19363
rect 10137 19323 10195 19329
rect 3602 19252 3608 19304
rect 3660 19292 3666 19304
rect 3786 19292 3792 19304
rect 3660 19264 3792 19292
rect 3660 19252 3666 19264
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 10060 19292 10088 19323
rect 9876 19264 10088 19292
rect 10152 19292 10180 19323
rect 10226 19320 10232 19372
rect 10284 19360 10290 19372
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 10284 19332 10329 19360
rect 10980 19332 12173 19360
rect 10284 19320 10290 19332
rect 10318 19292 10324 19304
rect 10152 19264 10324 19292
rect 9876 19236 9904 19264
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 10980 19292 11008 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12417 19363 12475 19369
rect 12417 19360 12429 19363
rect 12161 19323 12219 19329
rect 12268 19332 12429 19360
rect 10836 19264 11008 19292
rect 10836 19252 10842 19264
rect 11146 19252 11152 19304
rect 11204 19292 11210 19304
rect 12268 19292 12296 19332
rect 12417 19329 12429 19332
rect 12463 19329 12475 19363
rect 12417 19323 12475 19329
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19360 14795 19363
rect 16022 19360 16028 19372
rect 14783 19332 16028 19360
rect 14783 19329 14795 19332
rect 14737 19323 14795 19329
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 20714 19360 20720 19372
rect 20675 19332 20720 19360
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 21008 19369 21036 19400
rect 24026 19388 24032 19440
rect 24084 19428 24090 19440
rect 27264 19437 27292 19468
rect 30098 19456 30104 19468
rect 30156 19456 30162 19508
rect 27249 19431 27307 19437
rect 24084 19400 26096 19428
rect 24084 19388 24090 19400
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 21039 19332 22293 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 22462 19360 22468 19372
rect 22423 19332 22468 19360
rect 22281 19323 22339 19329
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 22925 19363 22983 19369
rect 22925 19329 22937 19363
rect 22971 19360 22983 19363
rect 23937 19363 23995 19369
rect 23937 19360 23949 19363
rect 22971 19332 23949 19360
rect 22971 19329 22983 19332
rect 22925 19323 22983 19329
rect 23937 19329 23949 19332
rect 23983 19329 23995 19363
rect 24118 19360 24124 19372
rect 24079 19332 24124 19360
rect 23937 19323 23995 19329
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24228 19369 24256 19400
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19329 24271 19363
rect 24486 19360 24492 19372
rect 24447 19332 24492 19360
rect 24213 19323 24271 19329
rect 24486 19320 24492 19332
rect 24544 19360 24550 19372
rect 25774 19360 25780 19372
rect 24544 19332 25780 19360
rect 24544 19320 24550 19332
rect 25774 19320 25780 19332
rect 25832 19320 25838 19372
rect 25958 19360 25964 19372
rect 25919 19332 25964 19360
rect 25958 19320 25964 19332
rect 26016 19320 26022 19372
rect 16942 19292 16948 19304
rect 11204 19264 12296 19292
rect 16903 19264 16948 19292
rect 11204 19252 11210 19264
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17218 19292 17224 19304
rect 17179 19264 17224 19292
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 20806 19292 20812 19304
rect 17328 19264 20668 19292
rect 20767 19264 20812 19292
rect 9858 19184 9864 19236
rect 9916 19184 9922 19236
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19224 14979 19227
rect 15010 19224 15016 19236
rect 14967 19196 15016 19224
rect 14967 19193 14979 19196
rect 14921 19187 14979 19193
rect 15010 19184 15016 19196
rect 15068 19224 15074 19236
rect 17328 19224 17356 19264
rect 15068 19196 17356 19224
rect 17681 19227 17739 19233
rect 15068 19184 15074 19196
rect 17681 19193 17693 19227
rect 17727 19224 17739 19227
rect 18046 19224 18052 19236
rect 17727 19196 18052 19224
rect 17727 19193 17739 19196
rect 17681 19187 17739 19193
rect 18046 19184 18052 19196
rect 18104 19184 18110 19236
rect 20533 19227 20591 19233
rect 20533 19224 20545 19227
rect 19904 19196 20545 19224
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 13446 19156 13452 19168
rect 10192 19128 13452 19156
rect 10192 19116 10198 19128
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 18690 19156 18696 19168
rect 13688 19128 18696 19156
rect 13688 19116 13694 19128
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19904 19165 19932 19196
rect 20533 19193 20545 19196
rect 20579 19193 20591 19227
rect 20640 19224 20668 19264
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 21174 19292 21180 19304
rect 20947 19264 21180 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 23198 19292 23204 19304
rect 23159 19264 23204 19292
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 23658 19252 23664 19304
rect 23716 19292 23722 19304
rect 24397 19295 24455 19301
rect 24397 19292 24409 19295
rect 23716 19264 24409 19292
rect 23716 19252 23722 19264
rect 24397 19261 24409 19264
rect 24443 19261 24455 19295
rect 24397 19255 24455 19261
rect 23750 19224 23756 19236
rect 20640 19196 23756 19224
rect 20533 19187 20591 19193
rect 23750 19184 23756 19196
rect 23808 19184 23814 19236
rect 26068 19224 26096 19400
rect 27249 19397 27261 19431
rect 27295 19397 27307 19431
rect 27249 19391 27307 19397
rect 28988 19431 29046 19437
rect 28988 19397 29000 19431
rect 29034 19428 29046 19431
rect 29822 19428 29828 19440
rect 29034 19400 29828 19428
rect 29034 19397 29046 19400
rect 28988 19391 29046 19397
rect 26145 19295 26203 19301
rect 26145 19261 26157 19295
rect 26191 19292 26203 19295
rect 27264 19292 27292 19391
rect 29822 19388 29828 19400
rect 29880 19388 29886 19440
rect 27614 19320 27620 19372
rect 27672 19360 27678 19372
rect 30561 19363 30619 19369
rect 27672 19332 30420 19360
rect 27672 19320 27678 19332
rect 26191 19264 27292 19292
rect 26191 19261 26203 19264
rect 26145 19255 26203 19261
rect 27982 19252 27988 19304
rect 28040 19292 28046 19304
rect 28721 19295 28779 19301
rect 28721 19292 28733 19295
rect 28040 19264 28733 19292
rect 28040 19252 28046 19264
rect 28721 19261 28733 19264
rect 28767 19261 28779 19295
rect 30392 19292 30420 19332
rect 30561 19329 30573 19363
rect 30607 19360 30619 19363
rect 30650 19360 30656 19372
rect 30607 19332 30656 19360
rect 30607 19329 30619 19332
rect 30561 19323 30619 19329
rect 30650 19320 30656 19332
rect 30708 19320 30714 19372
rect 30837 19295 30895 19301
rect 30837 19292 30849 19295
rect 30392 19264 30849 19292
rect 28721 19255 28779 19261
rect 30837 19261 30849 19264
rect 30883 19292 30895 19295
rect 30926 19292 30932 19304
rect 30883 19264 30932 19292
rect 30883 19261 30895 19264
rect 30837 19255 30895 19261
rect 30926 19252 30932 19264
rect 30984 19252 30990 19304
rect 26234 19224 26240 19236
rect 26068 19196 26240 19224
rect 26234 19184 26240 19196
rect 26292 19224 26298 19236
rect 27433 19227 27491 19233
rect 27433 19224 27445 19227
rect 26292 19196 27445 19224
rect 26292 19184 26298 19196
rect 27433 19193 27445 19196
rect 27479 19193 27491 19227
rect 27433 19187 27491 19193
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19125 19947 19159
rect 19889 19119 19947 19125
rect 22373 19159 22431 19165
rect 22373 19125 22385 19159
rect 22419 19156 22431 19159
rect 23017 19159 23075 19165
rect 23017 19156 23029 19159
rect 22419 19128 23029 19156
rect 22419 19125 22431 19128
rect 22373 19119 22431 19125
rect 23017 19125 23029 19128
rect 23063 19125 23075 19159
rect 23474 19156 23480 19168
rect 23435 19128 23480 19156
rect 23017 19119 23075 19125
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 27448 19156 27476 19187
rect 30466 19156 30472 19168
rect 27448 19128 30472 19156
rect 30466 19116 30472 19128
rect 30524 19116 30530 19168
rect 37829 19159 37887 19165
rect 37829 19125 37841 19159
rect 37875 19156 37887 19159
rect 38286 19156 38292 19168
rect 37875 19128 38292 19156
rect 37875 19125 37887 19128
rect 37829 19119 37887 19125
rect 38286 19116 38292 19128
rect 38344 19116 38350 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 9858 18952 9864 18964
rect 9447 18924 9864 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 10318 18952 10324 18964
rect 10279 18924 10324 18952
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 11974 18912 11980 18964
rect 12032 18952 12038 18964
rect 12161 18955 12219 18961
rect 12161 18952 12173 18955
rect 12032 18924 12173 18952
rect 12032 18912 12038 18924
rect 12161 18921 12173 18924
rect 12207 18921 12219 18955
rect 12161 18915 12219 18921
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 13504 18924 15240 18952
rect 13504 18912 13510 18924
rect 10686 18884 10692 18896
rect 4816 18856 10692 18884
rect 4816 18828 4844 18856
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 13541 18887 13599 18893
rect 13541 18884 13553 18887
rect 12406 18856 13553 18884
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 3326 18816 3332 18828
rect 2556 18788 3332 18816
rect 2556 18776 2562 18788
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 4798 18816 4804 18828
rect 4711 18788 4804 18816
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 8846 18776 8852 18828
rect 8904 18816 8910 18828
rect 10134 18816 10140 18828
rect 8904 18788 10140 18816
rect 8904 18776 8910 18788
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18748 2283 18751
rect 2777 18751 2835 18757
rect 2777 18748 2789 18751
rect 2271 18720 2789 18748
rect 2271 18717 2283 18720
rect 2225 18711 2283 18717
rect 2777 18717 2789 18720
rect 2823 18748 2835 18751
rect 9122 18748 9128 18760
rect 2823 18720 4016 18748
rect 9083 18720 9128 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 3988 18692 4016 18720
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9232 18757 9260 18788
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 10226 18748 10232 18760
rect 9539 18720 10232 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10778 18748 10784 18760
rect 10739 18720 10784 18748
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 11054 18757 11060 18760
rect 11048 18748 11060 18757
rect 11015 18720 11060 18748
rect 11048 18711 11060 18720
rect 11054 18708 11060 18711
rect 11112 18708 11118 18760
rect 2041 18683 2099 18689
rect 2041 18649 2053 18683
rect 2087 18680 2099 18683
rect 2958 18680 2964 18692
rect 2087 18652 2964 18680
rect 2087 18649 2099 18652
rect 2041 18643 2099 18649
rect 2240 18624 2268 18652
rect 2958 18640 2964 18652
rect 3016 18640 3022 18692
rect 3326 18680 3332 18692
rect 3287 18652 3332 18680
rect 3326 18640 3332 18652
rect 3384 18640 3390 18692
rect 3970 18680 3976 18692
rect 3931 18652 3976 18680
rect 3970 18640 3976 18652
rect 4028 18640 4034 18692
rect 9140 18680 9168 18708
rect 9140 18652 9444 18680
rect 2222 18572 2228 18624
rect 2280 18572 2286 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9416 18612 9444 18652
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 9953 18683 10011 18689
rect 9953 18680 9965 18683
rect 9640 18652 9965 18680
rect 9640 18640 9646 18652
rect 9953 18649 9965 18652
rect 9999 18680 10011 18683
rect 12406 18680 12434 18856
rect 13541 18853 13553 18856
rect 13587 18884 13599 18887
rect 13630 18884 13636 18896
rect 13587 18856 13636 18884
rect 13587 18853 13599 18856
rect 13541 18847 13599 18853
rect 13630 18844 13636 18856
rect 13688 18844 13694 18896
rect 15212 18884 15240 18924
rect 17218 18912 17224 18964
rect 17276 18952 17282 18964
rect 17773 18955 17831 18961
rect 17773 18952 17785 18955
rect 17276 18924 17785 18952
rect 17276 18912 17282 18924
rect 17773 18921 17785 18924
rect 17819 18921 17831 18955
rect 20162 18952 20168 18964
rect 20123 18924 20168 18952
rect 17773 18915 17831 18921
rect 20162 18912 20168 18924
rect 20220 18912 20226 18964
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 23477 18955 23535 18961
rect 23477 18952 23489 18955
rect 20864 18924 23489 18952
rect 20864 18912 20870 18924
rect 23477 18921 23489 18924
rect 23523 18921 23535 18955
rect 23477 18915 23535 18921
rect 31665 18955 31723 18961
rect 31665 18921 31677 18955
rect 31711 18952 31723 18955
rect 31846 18952 31852 18964
rect 31711 18924 31852 18952
rect 31711 18921 31723 18924
rect 31665 18915 31723 18921
rect 31846 18912 31852 18924
rect 31904 18912 31910 18964
rect 22370 18884 22376 18896
rect 15212 18856 22376 18884
rect 22370 18844 22376 18856
rect 22428 18844 22434 18896
rect 22462 18844 22468 18896
rect 22520 18884 22526 18896
rect 22925 18887 22983 18893
rect 22925 18884 22937 18887
rect 22520 18856 22937 18884
rect 22520 18844 22526 18856
rect 22925 18853 22937 18856
rect 22971 18853 22983 18887
rect 27430 18884 27436 18896
rect 27391 18856 27436 18884
rect 22925 18847 22983 18853
rect 27430 18844 27436 18856
rect 27488 18844 27494 18896
rect 28074 18844 28080 18896
rect 28132 18884 28138 18896
rect 28132 18856 28580 18884
rect 28132 18844 28138 18856
rect 17310 18816 17316 18828
rect 17271 18788 17316 18816
rect 17310 18776 17316 18788
rect 17368 18776 17374 18828
rect 20533 18819 20591 18825
rect 20533 18785 20545 18819
rect 20579 18816 20591 18819
rect 22738 18816 22744 18828
rect 20579 18788 22744 18816
rect 20579 18785 20591 18788
rect 20533 18779 20591 18785
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 25041 18819 25099 18825
rect 25041 18785 25053 18819
rect 25087 18816 25099 18819
rect 25958 18816 25964 18828
rect 25087 18788 25964 18816
rect 25087 18785 25099 18788
rect 25041 18779 25099 18785
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 28258 18816 28264 18828
rect 28219 18788 28264 18816
rect 28258 18776 28264 18788
rect 28316 18776 28322 18828
rect 28552 18760 28580 18856
rect 30650 18844 30656 18896
rect 30708 18884 30714 18896
rect 31021 18887 31079 18893
rect 31021 18884 31033 18887
rect 30708 18856 31033 18884
rect 30708 18844 30714 18856
rect 31021 18853 31033 18856
rect 31067 18853 31079 18887
rect 31021 18847 31079 18853
rect 31205 18819 31263 18825
rect 31205 18785 31217 18819
rect 31251 18816 31263 18819
rect 37826 18816 37832 18828
rect 31251 18788 31892 18816
rect 37787 18788 37832 18816
rect 31251 18785 31263 18788
rect 31205 18779 31263 18785
rect 13538 18708 13544 18760
rect 13596 18748 13602 18760
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13596 18720 13737 18748
rect 13596 18708 13602 18720
rect 13725 18717 13737 18720
rect 13771 18717 13783 18751
rect 13725 18711 13783 18717
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13872 18720 14289 18748
rect 13872 18708 13878 18720
rect 14277 18717 14289 18720
rect 14323 18717 14335 18751
rect 16117 18751 16175 18757
rect 16117 18748 16129 18751
rect 14277 18711 14335 18717
rect 15672 18720 16129 18748
rect 14550 18689 14556 18692
rect 9999 18652 12434 18680
rect 9999 18649 10011 18652
rect 9953 18643 10011 18649
rect 14544 18643 14556 18689
rect 14608 18680 14614 18692
rect 14608 18652 14644 18680
rect 14550 18640 14556 18643
rect 14608 18640 14614 18652
rect 10153 18615 10211 18621
rect 10153 18612 10165 18615
rect 9416 18584 10165 18612
rect 10153 18581 10165 18584
rect 10199 18581 10211 18615
rect 10153 18575 10211 18581
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 15672 18621 15700 18720
rect 16117 18717 16129 18720
rect 16163 18717 16175 18751
rect 16117 18711 16175 18717
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 16356 18720 17049 18748
rect 16356 18708 16362 18720
rect 17037 18717 17049 18720
rect 17083 18717 17095 18751
rect 17037 18711 17095 18717
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17405 18751 17463 18757
rect 17267 18720 17350 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17322 18624 17350 18720
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17600 18751 17658 18757
rect 17600 18717 17612 18751
rect 17646 18750 17658 18751
rect 17646 18748 17724 18750
rect 17646 18722 17816 18748
rect 17646 18717 17658 18722
rect 17696 18720 17816 18722
rect 17600 18711 17658 18717
rect 17420 18624 17448 18711
rect 15657 18615 15715 18621
rect 15657 18612 15669 18615
rect 15252 18584 15669 18612
rect 15252 18572 15258 18584
rect 15657 18581 15669 18584
rect 15703 18581 15715 18615
rect 15657 18575 15715 18581
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 15804 18584 16221 18612
rect 15804 18572 15810 18584
rect 16209 18581 16221 18584
rect 16255 18612 16267 18615
rect 17126 18612 17132 18624
rect 16255 18584 17132 18612
rect 16255 18581 16267 18584
rect 16209 18575 16267 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17310 18572 17316 18624
rect 17368 18572 17374 18624
rect 17402 18572 17408 18624
rect 17460 18572 17466 18624
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 17788 18612 17816 18720
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20441 18751 20499 18757
rect 20441 18748 20453 18751
rect 20404 18720 20453 18748
rect 20404 18708 20410 18720
rect 20441 18717 20453 18720
rect 20487 18717 20499 18751
rect 20622 18748 20628 18760
rect 20583 18720 20628 18748
rect 20441 18711 20499 18717
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21082 18748 21088 18760
rect 20947 18720 21088 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21082 18708 21088 18720
rect 21140 18708 21146 18760
rect 22186 18748 22192 18760
rect 22147 18720 22192 18748
rect 22186 18708 22192 18720
rect 22244 18708 22250 18760
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18748 23167 18751
rect 23198 18748 23204 18760
rect 23155 18720 23204 18748
rect 23155 18717 23167 18720
rect 23109 18711 23167 18717
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 24946 18748 24952 18760
rect 24907 18720 24952 18748
rect 24946 18708 24952 18720
rect 25004 18708 25010 18760
rect 27614 18748 27620 18760
rect 27575 18720 27620 18748
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 28442 18748 28448 18760
rect 28403 18720 28448 18748
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 31662 18748 31668 18760
rect 28592 18720 28685 18748
rect 31623 18720 31668 18748
rect 28592 18708 28598 18720
rect 31662 18708 31668 18720
rect 31720 18708 31726 18760
rect 31864 18757 31892 18788
rect 37826 18776 37832 18788
rect 37884 18776 37890 18828
rect 38102 18816 38108 18828
rect 38063 18788 38108 18816
rect 38102 18776 38108 18788
rect 38160 18776 38166 18828
rect 38286 18816 38292 18828
rect 38247 18788 38292 18816
rect 38286 18776 38292 18788
rect 38344 18776 38350 18828
rect 31849 18751 31907 18757
rect 31849 18717 31861 18751
rect 31895 18748 31907 18751
rect 32490 18748 32496 18760
rect 31895 18720 32496 18748
rect 31895 18717 31907 18720
rect 31849 18711 31907 18717
rect 32490 18708 32496 18720
rect 32548 18708 32554 18760
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 22370 18680 22376 18692
rect 17920 18652 22094 18680
rect 22331 18652 22376 18680
rect 17920 18640 17926 18652
rect 20806 18612 20812 18624
rect 17644 18584 17816 18612
rect 20767 18584 20812 18612
rect 17644 18572 17650 18584
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 22066 18612 22094 18652
rect 22370 18640 22376 18652
rect 22428 18640 22434 18692
rect 23842 18680 23848 18692
rect 22480 18652 23848 18680
rect 22480 18612 22508 18652
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 30466 18640 30472 18692
rect 30524 18680 30530 18692
rect 30745 18683 30803 18689
rect 30745 18680 30757 18683
rect 30524 18652 30757 18680
rect 30524 18640 30530 18652
rect 30745 18649 30757 18652
rect 30791 18649 30803 18683
rect 30745 18643 30803 18649
rect 23198 18612 23204 18624
rect 22066 18584 22508 18612
rect 23159 18584 23204 18612
rect 23198 18572 23204 18584
rect 23256 18572 23262 18624
rect 23293 18615 23351 18621
rect 23293 18581 23305 18615
rect 23339 18612 23351 18615
rect 24118 18612 24124 18624
rect 23339 18584 24124 18612
rect 23339 18581 23351 18584
rect 23293 18575 23351 18581
rect 24118 18572 24124 18584
rect 24176 18612 24182 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 24176 18584 24593 18612
rect 24176 18572 24182 18584
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 28258 18612 28264 18624
rect 28219 18584 28264 18612
rect 24581 18575 24639 18581
rect 28258 18572 28264 18584
rect 28316 18572 28322 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 11146 18408 11152 18420
rect 10459 18380 11152 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 12342 18408 12348 18420
rect 12303 18380 12348 18408
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 16114 18368 16120 18420
rect 16172 18408 16178 18420
rect 16853 18411 16911 18417
rect 16172 18380 16804 18408
rect 16172 18368 16178 18380
rect 4433 18343 4491 18349
rect 4433 18309 4445 18343
rect 4479 18340 4491 18343
rect 4614 18340 4620 18352
rect 4479 18312 4620 18340
rect 4479 18309 4491 18312
rect 4433 18303 4491 18309
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 9861 18343 9919 18349
rect 9861 18309 9873 18343
rect 9907 18340 9919 18343
rect 9907 18312 10548 18340
rect 9907 18309 9919 18312
rect 9861 18303 9919 18309
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4157 18275 4215 18281
rect 4157 18272 4169 18275
rect 4028 18244 4169 18272
rect 4028 18232 4034 18244
rect 4157 18241 4169 18244
rect 4203 18241 4215 18275
rect 8846 18272 8852 18284
rect 8807 18244 8852 18272
rect 4157 18235 4215 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18272 8999 18275
rect 9122 18272 9128 18284
rect 8987 18244 9128 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9582 18272 9588 18284
rect 9543 18244 9588 18272
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10318 18272 10324 18284
rect 10279 18244 10324 18272
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 10520 18281 10548 18312
rect 12158 18300 12164 18352
rect 12216 18340 12222 18352
rect 12989 18343 13047 18349
rect 12989 18340 13001 18343
rect 12216 18312 13001 18340
rect 12216 18300 12222 18312
rect 12989 18309 13001 18312
rect 13035 18309 13047 18343
rect 12989 18303 13047 18309
rect 14737 18343 14795 18349
rect 14737 18309 14749 18343
rect 14783 18340 14795 18343
rect 16574 18340 16580 18352
rect 14783 18312 16580 18340
rect 14783 18309 14795 18312
rect 14737 18303 14795 18309
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 16776 18340 16804 18380
rect 16853 18377 16865 18411
rect 16899 18408 16911 18411
rect 17678 18408 17684 18420
rect 16899 18380 17684 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 20622 18408 20628 18420
rect 20583 18380 20628 18408
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 22557 18411 22615 18417
rect 22557 18408 22569 18411
rect 22520 18380 22569 18408
rect 22520 18368 22526 18380
rect 22557 18377 22569 18380
rect 22603 18377 22615 18411
rect 22557 18371 22615 18377
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 23201 18411 23259 18417
rect 23201 18408 23213 18411
rect 22796 18380 23213 18408
rect 22796 18368 22802 18380
rect 23201 18377 23213 18380
rect 23247 18377 23259 18411
rect 28166 18408 28172 18420
rect 23201 18371 23259 18377
rect 27264 18380 28172 18408
rect 17218 18340 17224 18352
rect 16776 18312 17224 18340
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 18138 18340 18144 18352
rect 17512 18312 18144 18340
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18241 10563 18275
rect 10505 18235 10563 18241
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 11848 18244 12265 18272
rect 11848 18232 11854 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 12529 18275 12587 18281
rect 12529 18272 12541 18275
rect 12492 18244 12541 18272
rect 12492 18232 12498 18244
rect 12529 18241 12541 18244
rect 12575 18241 12587 18275
rect 15746 18272 15752 18284
rect 15707 18244 15752 18272
rect 12529 18235 12587 18241
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 1854 18204 1860 18216
rect 1815 18176 1860 18204
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 2038 18204 2044 18216
rect 1999 18176 2044 18204
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 2832 18176 2877 18204
rect 2832 18164 2838 18176
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9732 18176 9873 18204
rect 9732 18164 9738 18176
rect 9861 18173 9873 18176
rect 9907 18204 9919 18207
rect 15010 18204 15016 18216
rect 9907 18176 15016 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 16040 18204 16068 18235
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16172 18244 16217 18272
rect 16172 18232 16178 18244
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16356 18244 16401 18272
rect 16356 18232 16362 18244
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 16991 18275 17049 18281
rect 16991 18272 17003 18275
rect 16724 18244 17003 18272
rect 16724 18232 16730 18244
rect 16991 18241 17003 18244
rect 17037 18241 17049 18275
rect 17126 18272 17132 18284
rect 17087 18244 17132 18272
rect 16991 18235 17049 18241
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17512 18281 17540 18312
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 18693 18343 18751 18349
rect 18693 18340 18705 18343
rect 18472 18312 18705 18340
rect 18472 18300 18478 18312
rect 18693 18309 18705 18312
rect 18739 18309 18751 18343
rect 18693 18303 18751 18309
rect 20990 18300 20996 18352
rect 21048 18340 21054 18352
rect 25774 18340 25780 18352
rect 21048 18312 23428 18340
rect 25735 18312 25780 18340
rect 21048 18300 21054 18312
rect 17349 18275 17407 18281
rect 17349 18241 17361 18275
rect 17395 18241 17407 18275
rect 17349 18235 17407 18241
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 16758 18204 16764 18216
rect 16040 18176 16764 18204
rect 16758 18164 16764 18176
rect 16816 18204 16822 18216
rect 17364 18204 17392 18235
rect 17586 18232 17592 18284
rect 17644 18272 17650 18284
rect 20349 18275 20407 18281
rect 20349 18272 20361 18275
rect 17644 18244 20361 18272
rect 17644 18232 17650 18244
rect 20349 18241 20361 18244
rect 20395 18272 20407 18275
rect 20806 18272 20812 18284
rect 20395 18244 20812 18272
rect 20395 18241 20407 18244
rect 20349 18235 20407 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 23400 18281 23428 18312
rect 25774 18300 25780 18312
rect 25832 18300 25838 18352
rect 25866 18300 25872 18352
rect 25924 18340 25930 18352
rect 25961 18343 26019 18349
rect 25961 18340 25973 18343
rect 25924 18312 25973 18340
rect 25924 18300 25930 18312
rect 25961 18309 25973 18312
rect 26007 18340 26019 18343
rect 26050 18340 26056 18352
rect 26007 18312 26056 18340
rect 26007 18309 26019 18312
rect 25961 18303 26019 18309
rect 26050 18300 26056 18312
rect 26108 18300 26114 18352
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 23385 18275 23443 18281
rect 23385 18241 23397 18275
rect 23431 18241 23443 18275
rect 23385 18235 23443 18241
rect 16816 18176 17392 18204
rect 16816 18164 16822 18176
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 18288 18176 20637 18204
rect 18288 18164 18294 18176
rect 20625 18173 20637 18176
rect 20671 18204 20683 18207
rect 21174 18204 21180 18216
rect 20671 18176 21180 18204
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 21174 18164 21180 18176
rect 21232 18164 21238 18216
rect 15838 18136 15844 18148
rect 15799 18108 15844 18136
rect 15838 18096 15844 18108
rect 15896 18096 15902 18148
rect 17126 18096 17132 18148
rect 17184 18136 17190 18148
rect 17310 18136 17316 18148
rect 17184 18108 17316 18136
rect 17184 18096 17190 18108
rect 17310 18096 17316 18108
rect 17368 18136 17374 18148
rect 17368 18108 18368 18136
rect 17368 18096 17374 18108
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9677 18071 9735 18077
rect 9677 18068 9689 18071
rect 9171 18040 9689 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9677 18037 9689 18040
rect 9723 18068 9735 18071
rect 9858 18068 9864 18080
rect 9723 18040 9864 18068
rect 9723 18037 9735 18040
rect 9677 18031 9735 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 12529 18071 12587 18077
rect 12529 18037 12541 18071
rect 12575 18068 12587 18071
rect 12986 18068 12992 18080
rect 12575 18040 12992 18068
rect 12575 18037 12587 18040
rect 12529 18031 12587 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 13722 18028 13728 18080
rect 13780 18068 13786 18080
rect 17586 18068 17592 18080
rect 13780 18040 17592 18068
rect 13780 18028 13786 18040
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 18340 18068 18368 18108
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 22204 18136 22232 18235
rect 23474 18232 23480 18284
rect 23532 18272 23538 18284
rect 23658 18272 23664 18284
rect 23532 18244 23577 18272
rect 23619 18244 23664 18272
rect 23532 18232 23538 18244
rect 23658 18232 23664 18244
rect 23716 18232 23722 18284
rect 26510 18232 26516 18284
rect 26568 18272 26574 18284
rect 27264 18281 27292 18380
rect 28166 18368 28172 18380
rect 28224 18368 28230 18420
rect 31662 18408 31668 18420
rect 31623 18380 31668 18408
rect 31662 18368 31668 18380
rect 31720 18368 31726 18420
rect 30374 18300 30380 18352
rect 30432 18340 30438 18352
rect 30432 18312 30696 18340
rect 30432 18300 30438 18312
rect 27249 18275 27307 18281
rect 27249 18272 27261 18275
rect 26568 18244 27261 18272
rect 26568 18232 26574 18244
rect 27249 18241 27261 18244
rect 27295 18241 27307 18275
rect 27430 18272 27436 18284
rect 27391 18244 27436 18272
rect 27249 18235 27307 18241
rect 27430 18232 27436 18244
rect 27488 18232 27494 18284
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 27798 18272 27804 18284
rect 27571 18244 27804 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 27798 18232 27804 18244
rect 27856 18232 27862 18284
rect 27982 18272 27988 18284
rect 27943 18244 27988 18272
rect 27982 18232 27988 18244
rect 28040 18232 28046 18284
rect 28241 18275 28299 18281
rect 28241 18272 28253 18275
rect 28092 18244 28253 18272
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18204 22339 18207
rect 27154 18204 27160 18216
rect 22327 18176 27160 18204
rect 22327 18173 22339 18176
rect 22281 18167 22339 18173
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 28092 18204 28120 18244
rect 28241 18241 28253 18244
rect 28287 18241 28299 18275
rect 30466 18272 30472 18284
rect 28241 18235 28299 18241
rect 29380 18244 30472 18272
rect 27264 18176 28120 18204
rect 27264 18145 27292 18176
rect 18564 18108 22232 18136
rect 27249 18139 27307 18145
rect 18564 18096 18570 18108
rect 27249 18105 27261 18139
rect 27295 18105 27307 18139
rect 27249 18099 27307 18105
rect 18785 18071 18843 18077
rect 18785 18068 18797 18071
rect 18340 18040 18797 18068
rect 18785 18037 18797 18040
rect 18831 18037 18843 18071
rect 18785 18031 18843 18037
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 21082 18068 21088 18080
rect 20487 18040 21088 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 23566 18068 23572 18080
rect 23527 18040 23572 18068
rect 23566 18028 23572 18040
rect 23624 18028 23630 18080
rect 25958 18028 25964 18080
rect 26016 18068 26022 18080
rect 26145 18071 26203 18077
rect 26145 18068 26157 18071
rect 26016 18040 26157 18068
rect 26016 18028 26022 18040
rect 26145 18037 26157 18040
rect 26191 18037 26203 18071
rect 26145 18031 26203 18037
rect 27154 18028 27160 18080
rect 27212 18068 27218 18080
rect 29380 18077 29408 18244
rect 30466 18232 30472 18244
rect 30524 18232 30530 18284
rect 30668 18281 30696 18312
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18241 30711 18275
rect 30926 18272 30932 18284
rect 30887 18244 30932 18272
rect 30653 18235 30711 18241
rect 30926 18232 30932 18244
rect 30984 18232 30990 18284
rect 31478 18232 31484 18284
rect 31536 18272 31542 18284
rect 31573 18275 31631 18281
rect 31573 18272 31585 18275
rect 31536 18244 31585 18272
rect 31536 18232 31542 18244
rect 31573 18241 31585 18244
rect 31619 18241 31631 18275
rect 31573 18235 31631 18241
rect 31757 18275 31815 18281
rect 31757 18241 31769 18275
rect 31803 18272 31815 18275
rect 32030 18272 32036 18284
rect 31803 18244 32036 18272
rect 31803 18241 31815 18244
rect 31757 18235 31815 18241
rect 32030 18232 32036 18244
rect 32088 18272 32094 18284
rect 32309 18275 32367 18281
rect 32309 18272 32321 18275
rect 32088 18244 32321 18272
rect 32088 18232 32094 18244
rect 32309 18241 32321 18244
rect 32355 18241 32367 18275
rect 32490 18272 32496 18284
rect 32451 18244 32496 18272
rect 32309 18235 32367 18241
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 29365 18071 29423 18077
rect 29365 18068 29377 18071
rect 27212 18040 29377 18068
rect 27212 18028 27218 18040
rect 29365 18037 29377 18040
rect 29411 18037 29423 18071
rect 31110 18068 31116 18080
rect 31071 18040 31116 18068
rect 29365 18031 29423 18037
rect 31110 18028 31116 18040
rect 31168 18028 31174 18080
rect 31202 18028 31208 18080
rect 31260 18068 31266 18080
rect 32309 18071 32367 18077
rect 32309 18068 32321 18071
rect 31260 18040 32321 18068
rect 31260 18028 31266 18040
rect 32309 18037 32321 18040
rect 32355 18037 32367 18071
rect 32309 18031 32367 18037
rect 36446 18028 36452 18080
rect 36504 18068 36510 18080
rect 37461 18071 37519 18077
rect 37461 18068 37473 18071
rect 36504 18040 37473 18068
rect 36504 18028 36510 18040
rect 37461 18037 37473 18040
rect 37507 18037 37519 18071
rect 37461 18031 37519 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1765 17867 1823 17873
rect 1765 17833 1777 17867
rect 1811 17864 1823 17867
rect 1854 17864 1860 17876
rect 1811 17836 1860 17864
rect 1811 17833 1823 17836
rect 1765 17827 1823 17833
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2317 17867 2375 17873
rect 2317 17864 2329 17867
rect 2096 17836 2329 17864
rect 2096 17824 2102 17836
rect 2317 17833 2329 17836
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 9217 17867 9275 17873
rect 9217 17864 9229 17867
rect 9180 17836 9229 17864
rect 9180 17824 9186 17836
rect 9217 17833 9229 17836
rect 9263 17833 9275 17867
rect 13078 17864 13084 17876
rect 13039 17836 13084 17864
rect 9217 17827 9275 17833
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 14550 17864 14556 17876
rect 14511 17836 14556 17864
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 18138 17864 18144 17876
rect 18099 17836 18144 17864
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 23106 17864 23112 17876
rect 20180 17836 23112 17864
rect 9309 17799 9367 17805
rect 9309 17765 9321 17799
rect 9355 17796 9367 17799
rect 15562 17796 15568 17808
rect 9355 17768 9996 17796
rect 9355 17765 9367 17768
rect 9309 17759 9367 17765
rect 3602 17728 3608 17740
rect 2424 17700 3608 17728
rect 2424 17669 2452 17700
rect 3602 17688 3608 17700
rect 3660 17728 3666 17740
rect 4798 17728 4804 17740
rect 3660 17700 4804 17728
rect 3660 17688 3666 17700
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17728 9459 17731
rect 9674 17728 9680 17740
rect 9447 17700 9680 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 3234 17660 3240 17672
rect 3099 17632 3240 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 3970 17660 3976 17672
rect 3931 17632 3976 17660
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4706 17660 4712 17672
rect 4295 17632 4712 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8904 17632 9137 17660
rect 8904 17620 8910 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9858 17660 9864 17672
rect 9819 17632 9864 17660
rect 9125 17623 9183 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 9968 17660 9996 17768
rect 14844 17768 15568 17796
rect 10045 17663 10103 17669
rect 10045 17660 10057 17663
rect 9968 17632 10057 17660
rect 10045 17629 10057 17632
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 10778 17660 10784 17672
rect 10468 17632 10784 17660
rect 10468 17620 10474 17632
rect 10778 17620 10784 17632
rect 10836 17660 10842 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 10836 17632 11713 17660
rect 10836 17620 10842 17632
rect 11701 17629 11713 17632
rect 11747 17660 11759 17663
rect 13814 17660 13820 17672
rect 11747 17632 13820 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 14844 17669 14872 17768
rect 15562 17756 15568 17768
rect 15620 17756 15626 17808
rect 16206 17756 16212 17808
rect 16264 17796 16270 17808
rect 20180 17796 20208 17836
rect 23106 17824 23112 17836
rect 23164 17824 23170 17876
rect 27430 17824 27436 17876
rect 27488 17864 27494 17876
rect 27525 17867 27583 17873
rect 27525 17864 27537 17867
rect 27488 17836 27537 17864
rect 27488 17824 27494 17836
rect 27525 17833 27537 17836
rect 27571 17833 27583 17867
rect 27525 17827 27583 17833
rect 27798 17824 27804 17876
rect 27856 17864 27862 17876
rect 28077 17867 28135 17873
rect 28077 17864 28089 17867
rect 27856 17836 28089 17864
rect 27856 17824 27862 17836
rect 28077 17833 28089 17836
rect 28123 17833 28135 17867
rect 28077 17827 28135 17833
rect 30466 17824 30472 17876
rect 30524 17864 30530 17876
rect 32030 17864 32036 17876
rect 30524 17836 31892 17864
rect 31991 17836 32036 17864
rect 30524 17824 30530 17836
rect 20346 17796 20352 17808
rect 16264 17768 20208 17796
rect 20307 17768 20352 17796
rect 16264 17756 16270 17768
rect 20346 17756 20352 17768
rect 20404 17756 20410 17808
rect 28626 17796 28632 17808
rect 27632 17768 28632 17796
rect 16666 17728 16672 17740
rect 14936 17700 16672 17728
rect 14936 17669 14964 17700
rect 16666 17688 16672 17700
rect 16724 17728 16730 17740
rect 17310 17728 17316 17740
rect 16724 17700 17316 17728
rect 16724 17688 16730 17700
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17728 18659 17731
rect 19150 17728 19156 17740
rect 18647 17700 19156 17728
rect 18647 17697 18659 17700
rect 18601 17691 18659 17697
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 21174 17728 21180 17740
rect 20119 17700 21180 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 21174 17688 21180 17700
rect 21232 17688 21238 17740
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15010 17620 15016 17672
rect 15068 17660 15074 17672
rect 15194 17660 15200 17672
rect 15068 17632 15113 17660
rect 15155 17632 15200 17660
rect 15068 17620 15074 17632
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 18506 17660 18512 17672
rect 18467 17632 18512 17660
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 19978 17660 19984 17672
rect 19939 17632 19984 17660
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 25958 17660 25964 17672
rect 21048 17632 25452 17660
rect 25919 17632 25964 17660
rect 21048 17620 21054 17632
rect 9953 17595 10011 17601
rect 9953 17561 9965 17595
rect 9999 17592 10011 17595
rect 11946 17595 12004 17601
rect 11946 17592 11958 17595
rect 9999 17564 11958 17592
rect 9999 17561 10011 17564
rect 9953 17555 10011 17561
rect 11946 17561 11958 17564
rect 11992 17561 12004 17595
rect 13832 17592 13860 17620
rect 15657 17595 15715 17601
rect 15657 17592 15669 17595
rect 13832 17564 15669 17592
rect 11946 17555 12004 17561
rect 14936 17536 14964 17564
rect 15657 17561 15669 17564
rect 15703 17561 15715 17595
rect 15657 17555 15715 17561
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 17405 17595 17463 17601
rect 17405 17592 17417 17595
rect 16632 17564 17417 17592
rect 16632 17552 16638 17564
rect 17405 17561 17417 17564
rect 17451 17592 17463 17595
rect 22094 17592 22100 17604
rect 17451 17564 22100 17592
rect 17451 17561 17463 17564
rect 17405 17555 17463 17561
rect 22094 17552 22100 17564
rect 22152 17592 22158 17604
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 22152 17564 22569 17592
rect 22152 17552 22158 17564
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 22557 17555 22615 17561
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 24946 17592 24952 17604
rect 23072 17564 24952 17592
rect 23072 17552 23078 17564
rect 24946 17552 24952 17564
rect 25004 17552 25010 17604
rect 25424 17592 25452 17632
rect 25958 17620 25964 17632
rect 26016 17620 26022 17672
rect 26326 17660 26332 17672
rect 26287 17632 26332 17660
rect 26326 17620 26332 17632
rect 26384 17620 26390 17672
rect 26418 17620 26424 17672
rect 26476 17660 26482 17672
rect 26476 17632 26521 17660
rect 26476 17620 26482 17632
rect 27154 17620 27160 17672
rect 27212 17660 27218 17672
rect 27632 17669 27660 17768
rect 28626 17756 28632 17768
rect 28684 17796 28690 17808
rect 28994 17796 29000 17808
rect 28684 17768 29000 17796
rect 28684 17756 28690 17768
rect 28994 17756 29000 17768
rect 29052 17756 29058 17808
rect 31202 17796 31208 17808
rect 30852 17768 31208 17796
rect 30852 17737 30880 17768
rect 31202 17756 31208 17768
rect 31260 17756 31266 17808
rect 31864 17805 31892 17836
rect 32030 17824 32036 17836
rect 32088 17824 32094 17876
rect 31849 17799 31907 17805
rect 31849 17765 31861 17799
rect 31895 17765 31907 17799
rect 31849 17759 31907 17765
rect 30837 17731 30895 17737
rect 30837 17728 30849 17731
rect 28552 17700 30849 17728
rect 27433 17663 27491 17669
rect 27433 17660 27445 17663
rect 27212 17632 27445 17660
rect 27212 17620 27218 17632
rect 27433 17629 27445 17632
rect 27479 17629 27491 17663
rect 27433 17623 27491 17629
rect 27617 17663 27675 17669
rect 27617 17629 27629 17663
rect 27663 17629 27675 17663
rect 28258 17660 28264 17672
rect 28219 17632 28264 17660
rect 27617 17623 27675 17629
rect 28258 17620 28264 17632
rect 28316 17620 28322 17672
rect 28442 17620 28448 17672
rect 28500 17660 28506 17672
rect 28552 17669 28580 17700
rect 30837 17697 30849 17700
rect 30883 17697 30895 17731
rect 30837 17691 30895 17697
rect 31021 17731 31079 17737
rect 31021 17697 31033 17731
rect 31067 17728 31079 17731
rect 31110 17728 31116 17740
rect 31067 17700 31116 17728
rect 31067 17697 31079 17700
rect 31021 17691 31079 17697
rect 31110 17688 31116 17700
rect 31168 17688 31174 17740
rect 36446 17728 36452 17740
rect 36407 17700 36452 17728
rect 36446 17688 36452 17700
rect 36504 17688 36510 17740
rect 38286 17728 38292 17740
rect 38247 17700 38292 17728
rect 38286 17688 38292 17700
rect 38344 17688 38350 17740
rect 28537 17663 28595 17669
rect 28537 17660 28549 17663
rect 28500 17632 28549 17660
rect 28500 17620 28506 17632
rect 28537 17629 28549 17632
rect 28583 17629 28595 17663
rect 30742 17660 30748 17672
rect 30703 17632 30748 17660
rect 28537 17623 28595 17629
rect 30742 17620 30748 17632
rect 30800 17620 30806 17672
rect 30929 17663 30987 17669
rect 30929 17629 30941 17663
rect 30975 17660 30987 17663
rect 31478 17660 31484 17672
rect 30975 17632 31484 17660
rect 30975 17629 30987 17632
rect 30929 17623 30987 17629
rect 25682 17592 25688 17604
rect 25424 17564 25688 17592
rect 25682 17552 25688 17564
rect 25740 17592 25746 17604
rect 26053 17595 26111 17601
rect 26053 17592 26065 17595
rect 25740 17564 26065 17592
rect 25740 17552 25746 17564
rect 26053 17561 26065 17564
rect 26099 17561 26111 17595
rect 26053 17555 26111 17561
rect 2961 17527 3019 17533
rect 2961 17493 2973 17527
rect 3007 17524 3019 17527
rect 3510 17524 3516 17536
rect 3007 17496 3516 17524
rect 3007 17493 3019 17496
rect 2961 17487 3019 17493
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 14918 17484 14924 17536
rect 14976 17484 14982 17536
rect 16850 17484 16856 17536
rect 16908 17524 16914 17536
rect 17586 17524 17592 17536
rect 16908 17496 17592 17524
rect 16908 17484 16914 17496
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 22002 17524 22008 17536
rect 21315 17496 22008 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 23106 17484 23112 17536
rect 23164 17524 23170 17536
rect 25777 17527 25835 17533
rect 25777 17524 25789 17527
rect 23164 17496 25789 17524
rect 23164 17484 23170 17496
rect 25777 17493 25789 17496
rect 25823 17493 25835 17527
rect 26068 17524 26096 17555
rect 26142 17552 26148 17604
rect 26200 17592 26206 17604
rect 30944 17592 30972 17623
rect 31478 17620 31484 17632
rect 31536 17620 31542 17672
rect 26200 17564 26245 17592
rect 28552 17564 30972 17592
rect 26200 17552 26206 17564
rect 28552 17536 28580 17564
rect 31018 17552 31024 17604
rect 31076 17592 31082 17604
rect 31573 17595 31631 17601
rect 31573 17592 31585 17595
rect 31076 17564 31585 17592
rect 31076 17552 31082 17564
rect 31573 17561 31585 17564
rect 31619 17561 31631 17595
rect 31573 17555 31631 17561
rect 36633 17595 36691 17601
rect 36633 17561 36645 17595
rect 36679 17592 36691 17595
rect 37550 17592 37556 17604
rect 36679 17564 37556 17592
rect 36679 17561 36691 17564
rect 36633 17555 36691 17561
rect 37550 17552 37556 17564
rect 37608 17552 37614 17604
rect 27154 17524 27160 17536
rect 26068 17496 27160 17524
rect 25777 17487 25835 17493
rect 27154 17484 27160 17496
rect 27212 17484 27218 17536
rect 28445 17527 28503 17533
rect 28445 17493 28457 17527
rect 28491 17524 28503 17527
rect 28534 17524 28540 17536
rect 28491 17496 28540 17524
rect 28491 17493 28503 17496
rect 28445 17487 28503 17493
rect 28534 17484 28540 17496
rect 28592 17484 28598 17536
rect 30282 17484 30288 17536
rect 30340 17524 30346 17536
rect 30561 17527 30619 17533
rect 30561 17524 30573 17527
rect 30340 17496 30573 17524
rect 30340 17484 30346 17496
rect 30561 17493 30573 17496
rect 30607 17493 30619 17527
rect 30561 17487 30619 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 3234 17280 3240 17332
rect 3292 17320 3298 17332
rect 3292 17292 22324 17320
rect 3292 17280 3298 17292
rect 3510 17252 3516 17264
rect 3471 17224 3516 17252
rect 3510 17212 3516 17224
rect 3568 17212 3574 17264
rect 12618 17212 12624 17264
rect 12676 17252 12682 17264
rect 13538 17252 13544 17264
rect 12676 17224 13544 17252
rect 12676 17212 12682 17224
rect 13538 17212 13544 17224
rect 13596 17252 13602 17264
rect 16942 17252 16948 17264
rect 13596 17224 16948 17252
rect 13596 17212 13602 17224
rect 16942 17212 16948 17224
rect 17000 17212 17006 17264
rect 17310 17252 17316 17264
rect 17271 17224 17316 17252
rect 17310 17212 17316 17224
rect 17368 17212 17374 17264
rect 17681 17255 17739 17261
rect 17681 17221 17693 17255
rect 17727 17252 17739 17255
rect 17770 17252 17776 17264
rect 17727 17224 17776 17252
rect 17727 17221 17739 17224
rect 17681 17215 17739 17221
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 21082 17252 21088 17264
rect 21043 17224 21088 17252
rect 21082 17212 21088 17224
rect 21140 17212 21146 17264
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 13630 17184 13636 17196
rect 13311 17156 13636 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 13814 17184 13820 17196
rect 13775 17156 13820 17184
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14084 17187 14142 17193
rect 14084 17153 14096 17187
rect 14130 17184 14142 17187
rect 14642 17184 14648 17196
rect 14130 17156 14648 17184
rect 14130 17153 14142 17156
rect 14084 17147 14142 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 16022 17144 16028 17196
rect 16080 17193 16086 17196
rect 16080 17187 16108 17193
rect 16096 17184 16108 17187
rect 17494 17184 17500 17196
rect 16096 17156 17172 17184
rect 17455 17156 17500 17184
rect 16096 17153 16108 17156
rect 16080 17147 16108 17153
rect 16080 17144 16086 17147
rect 1854 17116 1860 17128
rect 1815 17088 1860 17116
rect 1854 17076 1860 17088
rect 1912 17076 1918 17128
rect 2130 17076 2136 17128
rect 2188 17116 2194 17128
rect 3697 17119 3755 17125
rect 3697 17116 3709 17119
rect 2188 17088 3709 17116
rect 2188 17076 2194 17088
rect 3697 17085 3709 17088
rect 3743 17085 3755 17119
rect 17144 17116 17172 17156
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 19426 17184 19432 17196
rect 19387 17156 19432 17184
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20990 17184 20996 17196
rect 19536 17156 20996 17184
rect 19334 17116 19340 17128
rect 17144 17088 19340 17116
rect 3697 17079 3755 17085
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 19536 17125 19564 17156
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 21174 17184 21180 17196
rect 21135 17156 21180 17184
rect 21174 17144 21180 17156
rect 21232 17184 21238 17196
rect 21232 17156 22094 17184
rect 21232 17144 21238 17156
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 12894 17008 12900 17060
rect 12952 17048 12958 17060
rect 13081 17051 13139 17057
rect 13081 17048 13093 17051
rect 12952 17020 13093 17048
rect 12952 17008 12958 17020
rect 13081 17017 13093 17020
rect 13127 17017 13139 17051
rect 13081 17011 13139 17017
rect 13170 17008 13176 17060
rect 13228 17048 13234 17060
rect 15197 17051 15255 17057
rect 13228 17020 13273 17048
rect 13228 17008 13234 17020
rect 15197 17017 15209 17051
rect 15243 17048 15255 17051
rect 17034 17048 17040 17060
rect 15243 17020 17040 17048
rect 15243 17017 15255 17020
rect 15197 17011 15255 17017
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 14182 16980 14188 16992
rect 12851 16952 14188 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 15212 16980 15240 17011
rect 17034 17008 17040 17020
rect 17092 17008 17098 17060
rect 19797 17051 19855 17057
rect 19797 17017 19809 17051
rect 19843 17048 19855 17051
rect 19978 17048 19984 17060
rect 19843 17020 19984 17048
rect 19843 17017 19855 17020
rect 19797 17011 19855 17017
rect 19978 17008 19984 17020
rect 20036 17008 20042 17060
rect 22066 17048 22094 17156
rect 22296 17116 22324 17292
rect 23198 17280 23204 17332
rect 23256 17280 23262 17332
rect 23658 17280 23664 17332
rect 23716 17320 23722 17332
rect 23937 17323 23995 17329
rect 23937 17320 23949 17323
rect 23716 17292 23949 17320
rect 23716 17280 23722 17292
rect 23937 17289 23949 17292
rect 23983 17289 23995 17323
rect 23937 17283 23995 17289
rect 25945 17323 26003 17329
rect 25945 17289 25957 17323
rect 25991 17320 26003 17323
rect 26050 17320 26056 17332
rect 25991 17292 26056 17320
rect 25991 17289 26003 17292
rect 25945 17283 26003 17289
rect 26050 17280 26056 17292
rect 26108 17320 26114 17332
rect 26108 17292 26280 17320
rect 26108 17280 26114 17292
rect 23106 17252 23112 17264
rect 23067 17224 23112 17252
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 23216 17252 23244 17280
rect 26145 17255 26203 17261
rect 23216 17224 24348 17252
rect 22370 17144 22376 17196
rect 22428 17184 22434 17196
rect 22925 17187 22983 17193
rect 22925 17184 22937 17187
rect 22428 17156 22937 17184
rect 22428 17144 22434 17156
rect 22925 17153 22937 17156
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 23014 17144 23020 17196
rect 23072 17184 23078 17196
rect 23201 17187 23259 17193
rect 23201 17184 23213 17187
rect 23072 17156 23213 17184
rect 23072 17144 23078 17156
rect 23201 17153 23213 17156
rect 23247 17153 23259 17187
rect 23201 17147 23259 17153
rect 23290 17144 23296 17196
rect 23348 17184 23354 17196
rect 24320 17193 24348 17224
rect 26145 17221 26157 17255
rect 26191 17221 26203 17255
rect 26252 17252 26280 17292
rect 26326 17280 26332 17332
rect 26384 17320 26390 17332
rect 27249 17323 27307 17329
rect 27249 17320 27261 17323
rect 26384 17292 27261 17320
rect 26384 17280 26390 17292
rect 27249 17289 27261 17292
rect 27295 17289 27307 17323
rect 30282 17320 30288 17332
rect 30243 17292 30288 17320
rect 27249 17283 27307 17289
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 37550 17320 37556 17332
rect 37511 17292 37556 17320
rect 37550 17280 37556 17292
rect 37608 17280 37614 17332
rect 26252 17224 27476 17252
rect 26145 17215 26203 17221
rect 24305 17187 24363 17193
rect 23348 17156 23393 17184
rect 23492 17156 24164 17184
rect 23348 17144 23354 17156
rect 23382 17116 23388 17128
rect 22296 17088 23388 17116
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 23492 17048 23520 17156
rect 22066 17020 23520 17048
rect 23566 17008 23572 17060
rect 23624 17048 23630 17060
rect 24136 17048 24164 17156
rect 24305 17153 24317 17187
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 25133 17187 25191 17193
rect 25133 17153 25145 17187
rect 25179 17153 25191 17187
rect 25133 17147 25191 17153
rect 24397 17119 24455 17125
rect 24397 17085 24409 17119
rect 24443 17116 24455 17119
rect 25148 17116 25176 17147
rect 24443 17088 25176 17116
rect 24443 17085 24455 17088
rect 24397 17079 24455 17085
rect 24949 17051 25007 17057
rect 24949 17048 24961 17051
rect 23624 17020 23888 17048
rect 24136 17020 24961 17048
rect 23624 17008 23630 17020
rect 14516 16952 15240 16980
rect 14516 16940 14522 16952
rect 15286 16940 15292 16992
rect 15344 16980 15350 16992
rect 16206 16980 16212 16992
rect 15344 16952 16212 16980
rect 15344 16940 15350 16952
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 17954 16980 17960 16992
rect 17000 16952 17960 16980
rect 17000 16940 17006 16952
rect 17954 16940 17960 16952
rect 18012 16980 18018 16992
rect 23014 16980 23020 16992
rect 18012 16952 23020 16980
rect 18012 16940 18018 16952
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 23477 16983 23535 16989
rect 23477 16949 23489 16983
rect 23523 16980 23535 16983
rect 23750 16980 23756 16992
rect 23523 16952 23756 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 23750 16940 23756 16952
rect 23808 16940 23814 16992
rect 23860 16980 23888 17020
rect 24949 17017 24961 17020
rect 24995 17017 25007 17051
rect 25148 17048 25176 17088
rect 25314 17076 25320 17128
rect 25372 17116 25378 17128
rect 26050 17116 26056 17128
rect 25372 17088 26056 17116
rect 25372 17076 25378 17088
rect 26050 17076 26056 17088
rect 26108 17076 26114 17128
rect 26160 17116 26188 17215
rect 27448 17196 27476 17224
rect 27154 17184 27160 17196
rect 27115 17156 27160 17184
rect 27154 17144 27160 17156
rect 27212 17144 27218 17196
rect 27430 17184 27436 17196
rect 27343 17156 27436 17184
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 30098 17184 30104 17196
rect 30059 17156 30104 17184
rect 30098 17144 30104 17156
rect 30156 17144 30162 17196
rect 30374 17144 30380 17196
rect 30432 17184 30438 17196
rect 36909 17187 36967 17193
rect 30432 17156 30477 17184
rect 30432 17144 30438 17156
rect 36909 17153 36921 17187
rect 36955 17184 36967 17187
rect 37274 17184 37280 17196
rect 36955 17156 37280 17184
rect 36955 17153 36967 17156
rect 36909 17147 36967 17153
rect 37274 17144 37280 17156
rect 37332 17144 37338 17196
rect 37645 17187 37703 17193
rect 37645 17153 37657 17187
rect 37691 17184 37703 17187
rect 38010 17184 38016 17196
rect 37691 17156 38016 17184
rect 37691 17153 37703 17156
rect 37645 17147 37703 17153
rect 38010 17144 38016 17156
rect 38068 17144 38074 17196
rect 26234 17116 26240 17128
rect 26160 17088 26240 17116
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 27525 17119 27583 17125
rect 27525 17085 27537 17119
rect 27571 17116 27583 17119
rect 27614 17116 27620 17128
rect 27571 17088 27620 17116
rect 27571 17085 27583 17088
rect 27525 17079 27583 17085
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 25777 17051 25835 17057
rect 25777 17048 25789 17051
rect 25148 17020 25789 17048
rect 24949 17011 25007 17017
rect 25777 17017 25789 17020
rect 25823 17017 25835 17051
rect 33870 17048 33876 17060
rect 25777 17011 25835 17017
rect 25884 17020 33876 17048
rect 25884 16980 25912 17020
rect 33870 17008 33876 17020
rect 33928 17008 33934 17060
rect 23860 16952 25912 16980
rect 25958 16940 25964 16992
rect 26016 16980 26022 16992
rect 26016 16952 26061 16980
rect 26016 16940 26022 16952
rect 26142 16940 26148 16992
rect 26200 16980 26206 16992
rect 27338 16980 27344 16992
rect 26200 16952 27344 16980
rect 26200 16940 26206 16952
rect 27338 16940 27344 16952
rect 27396 16940 27402 16992
rect 28350 16940 28356 16992
rect 28408 16980 28414 16992
rect 30101 16983 30159 16989
rect 30101 16980 30113 16983
rect 28408 16952 30113 16980
rect 28408 16940 28414 16952
rect 30101 16949 30113 16952
rect 30147 16949 30159 16983
rect 30101 16943 30159 16949
rect 36630 16940 36636 16992
rect 36688 16980 36694 16992
rect 36817 16983 36875 16989
rect 36817 16980 36829 16983
rect 36688 16952 36829 16980
rect 36688 16940 36694 16952
rect 36817 16949 36829 16952
rect 36863 16949 36875 16983
rect 38102 16980 38108 16992
rect 38063 16952 38108 16980
rect 36817 16943 36875 16949
rect 38102 16940 38108 16952
rect 38160 16940 38166 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2130 16776 2136 16788
rect 2091 16748 2136 16776
rect 2130 16736 2136 16748
rect 2188 16736 2194 16788
rect 3786 16736 3792 16788
rect 3844 16776 3850 16788
rect 3970 16776 3976 16788
rect 3844 16748 3976 16776
rect 3844 16736 3850 16748
rect 3970 16736 3976 16748
rect 4028 16776 4034 16788
rect 12894 16776 12900 16788
rect 4028 16748 12756 16776
rect 12855 16748 12900 16776
rect 4028 16736 4034 16748
rect 10781 16711 10839 16717
rect 10781 16677 10793 16711
rect 10827 16708 10839 16711
rect 12618 16708 12624 16720
rect 10827 16680 11192 16708
rect 10827 16677 10839 16680
rect 10781 16671 10839 16677
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 9217 16643 9275 16649
rect 9217 16640 9229 16643
rect 9180 16612 9229 16640
rect 9180 16600 9186 16612
rect 9217 16609 9229 16612
rect 9263 16609 9275 16643
rect 10502 16640 10508 16652
rect 10463 16612 10508 16640
rect 9217 16603 9275 16609
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 4430 16572 4436 16584
rect 3467 16544 4436 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 9309 16575 9367 16581
rect 9309 16572 9321 16575
rect 8904 16544 9321 16572
rect 8904 16532 8910 16544
rect 9309 16541 9321 16544
rect 9355 16541 9367 16575
rect 9309 16535 9367 16541
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 10284 16544 10425 16572
rect 10284 16532 10290 16544
rect 10413 16541 10425 16544
rect 10459 16541 10471 16575
rect 11164 16572 11192 16680
rect 11624 16680 12624 16708
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11624 16640 11652 16680
rect 12618 16668 12624 16680
rect 12676 16668 12682 16720
rect 12728 16708 12756 16748
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 13228 16748 13461 16776
rect 13228 16736 13234 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 13630 16736 13636 16788
rect 13688 16776 13694 16788
rect 14458 16776 14464 16788
rect 13688 16748 14464 16776
rect 13688 16736 13694 16748
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 14737 16779 14795 16785
rect 14737 16776 14749 16779
rect 14700 16748 14749 16776
rect 14700 16736 14706 16748
rect 14737 16745 14749 16748
rect 14783 16745 14795 16779
rect 14737 16739 14795 16745
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 16853 16779 16911 16785
rect 16853 16776 16865 16779
rect 16816 16748 16865 16776
rect 16816 16736 16822 16748
rect 16853 16745 16865 16748
rect 16899 16745 16911 16779
rect 16853 16739 16911 16745
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 17678 16776 17684 16788
rect 17460 16748 17684 16776
rect 17460 16736 17466 16748
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 20993 16779 21051 16785
rect 20993 16745 21005 16779
rect 21039 16776 21051 16779
rect 21637 16779 21695 16785
rect 21637 16776 21649 16779
rect 21039 16748 21649 16776
rect 21039 16745 21051 16748
rect 20993 16739 21051 16745
rect 21637 16745 21649 16748
rect 21683 16745 21695 16779
rect 21637 16739 21695 16745
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 27672 16748 30328 16776
rect 27672 16736 27678 16748
rect 30300 16717 30328 16748
rect 30374 16736 30380 16788
rect 30432 16776 30438 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 30432 16748 31217 16776
rect 30432 16736 30438 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 38010 16776 38016 16788
rect 31205 16739 31263 16745
rect 35866 16748 38016 16776
rect 30285 16711 30343 16717
rect 12728 16680 28488 16708
rect 11287 16612 11652 16640
rect 11793 16643 11851 16649
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 11839 16612 14136 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 12434 16581 12440 16584
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 11164 16544 11529 16572
rect 10413 16535 10471 16541
rect 11517 16541 11529 16544
rect 11563 16541 11575 16575
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11517 16535 11575 16541
rect 11624 16544 12265 16572
rect 3145 16507 3203 16513
rect 3145 16473 3157 16507
rect 3191 16473 3203 16507
rect 3145 16467 3203 16473
rect 4157 16507 4215 16513
rect 4157 16473 4169 16507
rect 4203 16504 4215 16507
rect 4798 16504 4804 16516
rect 4203 16476 4804 16504
rect 4203 16473 4215 16476
rect 4157 16467 4215 16473
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3160 16436 3188 16467
rect 4798 16464 4804 16476
rect 4856 16464 4862 16516
rect 11624 16513 11652 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12391 16575 12440 16581
rect 12391 16572 12403 16575
rect 12347 16544 12403 16572
rect 12253 16535 12311 16541
rect 12391 16541 12403 16544
rect 12437 16541 12440 16575
rect 12391 16535 12440 16541
rect 12434 16532 12440 16535
rect 12492 16532 12498 16584
rect 12718 16575 12776 16581
rect 12718 16541 12730 16575
rect 12764 16572 12776 16575
rect 13354 16572 13360 16584
rect 12764 16544 12848 16572
rect 13315 16544 13360 16572
rect 12764 16541 12776 16544
rect 12718 16535 12776 16541
rect 11609 16507 11667 16513
rect 11609 16504 11621 16507
rect 9692 16476 11621 16504
rect 8478 16436 8484 16448
rect 3016 16408 8484 16436
rect 3016 16396 3022 16408
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 9692 16445 9720 16476
rect 11609 16473 11621 16476
rect 11655 16473 11667 16507
rect 11609 16467 11667 16473
rect 11790 16464 11796 16516
rect 11848 16504 11854 16516
rect 12529 16507 12587 16513
rect 12529 16504 12541 16507
rect 11848 16476 12541 16504
rect 11848 16464 11854 16476
rect 12529 16473 12541 16476
rect 12575 16473 12587 16507
rect 12529 16467 12587 16473
rect 12618 16464 12624 16516
rect 12676 16504 12682 16516
rect 12676 16476 12721 16504
rect 12676 16464 12682 16476
rect 9677 16439 9735 16445
rect 9677 16405 9689 16439
rect 9723 16405 9735 16439
rect 11422 16436 11428 16448
rect 11383 16408 11428 16436
rect 9677 16399 9735 16405
rect 11422 16396 11428 16408
rect 11480 16436 11486 16448
rect 12820 16436 12848 16544
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13538 16572 13544 16584
rect 13499 16544 13544 16572
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 14108 16572 14136 16612
rect 14182 16600 14188 16652
rect 14240 16640 14246 16652
rect 14277 16643 14335 16649
rect 14277 16640 14289 16643
rect 14240 16612 14289 16640
rect 14240 16600 14246 16612
rect 14277 16609 14289 16612
rect 14323 16609 14335 16643
rect 16850 16640 16856 16652
rect 14277 16603 14335 16609
rect 15856 16612 16856 16640
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 14108 16544 14381 16572
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 15286 16572 15292 16584
rect 14599 16544 15292 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 14384 16504 14412 16535
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 15856 16581 15884 16612
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 25777 16643 25835 16649
rect 25777 16609 25789 16643
rect 25823 16640 25835 16643
rect 25866 16640 25872 16652
rect 25823 16612 25872 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 25866 16600 25872 16612
rect 25924 16600 25930 16652
rect 25958 16600 25964 16652
rect 26016 16640 26022 16652
rect 26053 16643 26111 16649
rect 26053 16640 26065 16643
rect 26016 16612 26065 16640
rect 26016 16600 26022 16612
rect 26053 16609 26065 16612
rect 26099 16640 26111 16643
rect 27614 16640 27620 16652
rect 26099 16612 27620 16640
rect 26099 16609 26111 16612
rect 26053 16603 26111 16609
rect 27614 16600 27620 16612
rect 27672 16600 27678 16652
rect 28350 16640 28356 16652
rect 28311 16612 28356 16640
rect 28350 16600 28356 16612
rect 28408 16600 28414 16652
rect 28460 16640 28488 16680
rect 30285 16677 30297 16711
rect 30331 16708 30343 16711
rect 30466 16708 30472 16720
rect 30331 16680 30472 16708
rect 30331 16677 30343 16680
rect 30285 16671 30343 16677
rect 30466 16668 30472 16680
rect 30524 16668 30530 16720
rect 35866 16640 35894 16748
rect 38010 16736 38016 16748
rect 38068 16736 38074 16788
rect 38102 16708 38108 16720
rect 36464 16680 38108 16708
rect 36464 16649 36492 16680
rect 38102 16668 38108 16680
rect 38160 16668 38166 16720
rect 28460 16612 35894 16640
rect 36449 16643 36507 16649
rect 36449 16609 36461 16643
rect 36495 16609 36507 16643
rect 36630 16640 36636 16652
rect 36591 16612 36636 16640
rect 36449 16603 36507 16609
rect 36630 16600 36636 16612
rect 36688 16600 36694 16652
rect 38286 16640 38292 16652
rect 38247 16612 38292 16640
rect 38286 16600 38292 16612
rect 38344 16600 38350 16652
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 15841 16535 15899 16541
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16942 16572 16948 16584
rect 16903 16544 16948 16572
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17586 16572 17592 16584
rect 17547 16544 17592 16572
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 18233 16575 18291 16581
rect 17736 16566 18184 16572
rect 18233 16566 18245 16575
rect 17736 16544 18245 16566
rect 17736 16532 17742 16544
rect 18156 16541 18245 16544
rect 18279 16541 18291 16575
rect 18156 16538 18291 16541
rect 18233 16535 18291 16538
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 18506 16572 18512 16584
rect 18463 16544 18512 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20640 16504 20668 16535
rect 21726 16532 21732 16584
rect 21784 16572 21790 16584
rect 21821 16575 21879 16581
rect 21821 16572 21833 16575
rect 21784 16544 21833 16572
rect 21784 16532 21790 16544
rect 21821 16541 21833 16544
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16572 22155 16575
rect 23290 16572 23296 16584
rect 22143 16544 23296 16572
rect 22143 16541 22155 16544
rect 22097 16535 22155 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 28258 16572 28264 16584
rect 28219 16544 28264 16572
rect 28258 16532 28264 16544
rect 28316 16532 28322 16584
rect 30653 16575 30711 16581
rect 30653 16541 30665 16575
rect 30699 16572 30711 16575
rect 30926 16572 30932 16584
rect 30699 16544 30932 16572
rect 30699 16541 30711 16544
rect 30653 16535 30711 16541
rect 30926 16532 30932 16544
rect 30984 16532 30990 16584
rect 31294 16572 31300 16584
rect 31255 16544 31300 16572
rect 31294 16532 31300 16544
rect 31352 16532 31358 16584
rect 14384 16476 15792 16504
rect 15654 16436 15660 16448
rect 11480 16408 12848 16436
rect 15615 16408 15660 16436
rect 11480 16396 11486 16408
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 15764 16436 15792 16476
rect 16960 16476 20668 16504
rect 16960 16436 16988 16476
rect 18230 16436 18236 16448
rect 15764 16408 16988 16436
rect 18191 16408 18236 16436
rect 18230 16396 18236 16408
rect 18288 16396 18294 16448
rect 20990 16436 20996 16448
rect 20951 16408 20996 16436
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 21177 16439 21235 16445
rect 21177 16405 21189 16439
rect 21223 16436 21235 16439
rect 21266 16436 21272 16448
rect 21223 16408 21272 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 21818 16396 21824 16448
rect 21876 16436 21882 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21876 16408 22017 16436
rect 21876 16396 21882 16408
rect 22005 16405 22017 16408
rect 22051 16436 22063 16439
rect 23750 16436 23756 16448
rect 22051 16408 23756 16436
rect 22051 16405 22063 16408
rect 22005 16399 22063 16405
rect 23750 16396 23756 16408
rect 23808 16436 23814 16448
rect 24302 16436 24308 16448
rect 23808 16408 24308 16436
rect 23808 16396 23814 16408
rect 24302 16396 24308 16408
rect 24360 16396 24366 16448
rect 27890 16436 27896 16448
rect 27851 16408 27896 16436
rect 27890 16396 27896 16408
rect 27948 16396 27954 16448
rect 30098 16396 30104 16448
rect 30156 16436 30162 16448
rect 30193 16439 30251 16445
rect 30193 16436 30205 16439
rect 30156 16408 30205 16436
rect 30156 16396 30162 16408
rect 30193 16405 30205 16408
rect 30239 16405 30251 16439
rect 30193 16399 30251 16405
rect 30282 16396 30288 16448
rect 30340 16436 30346 16448
rect 37366 16436 37372 16448
rect 30340 16408 37372 16436
rect 30340 16396 30346 16408
rect 37366 16396 37372 16408
rect 37424 16396 37430 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12802 16232 12808 16244
rect 12492 16204 12808 16232
rect 12492 16192 12498 16204
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 16850 16232 16856 16244
rect 16811 16204 16856 16232
rect 16850 16192 16856 16204
rect 16908 16192 16914 16244
rect 17218 16232 17224 16244
rect 17144 16204 17224 16232
rect 3145 16167 3203 16173
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 3234 16164 3240 16176
rect 3191 16136 3240 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 3694 16124 3700 16176
rect 3752 16164 3758 16176
rect 17144 16173 17172 16204
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 23290 16192 23296 16244
rect 23348 16232 23354 16244
rect 23385 16235 23443 16241
rect 23385 16232 23397 16235
rect 23348 16204 23397 16232
rect 23348 16192 23354 16204
rect 23385 16201 23397 16204
rect 23431 16201 23443 16235
rect 23385 16195 23443 16201
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 3752 16136 4537 16164
rect 3752 16124 3758 16136
rect 4525 16133 4537 16136
rect 4571 16164 4583 16167
rect 17129 16167 17187 16173
rect 4571 16136 12434 16164
rect 4571 16133 4583 16136
rect 4525 16127 4583 16133
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 2455 16068 2881 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2869 16065 2881 16068
rect 2915 16096 2927 16099
rect 3789 16099 3847 16105
rect 3789 16096 3801 16099
rect 2915 16068 3801 16096
rect 2915 16065 2927 16068
rect 2869 16059 2927 16065
rect 3789 16065 3801 16068
rect 3835 16096 3847 16099
rect 4430 16096 4436 16108
rect 3835 16068 4436 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4430 16056 4436 16068
rect 4488 16096 4494 16108
rect 4614 16096 4620 16108
rect 4488 16068 4620 16096
rect 4488 16056 4494 16068
rect 4614 16056 4620 16068
rect 4672 16096 4678 16108
rect 5261 16099 5319 16105
rect 5261 16096 5273 16099
rect 4672 16068 5273 16096
rect 4672 16056 4678 16068
rect 5261 16065 5273 16068
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 10284 16068 10425 16096
rect 10284 16056 10290 16068
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 15997 5871 16031
rect 10502 16028 10508 16040
rect 10463 16000 10508 16028
rect 5813 15991 5871 15997
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 5828 15960 5856 15991
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 10781 16031 10839 16037
rect 10781 15997 10793 16031
rect 10827 16028 10839 16031
rect 11790 16028 11796 16040
rect 10827 16000 11796 16028
rect 10827 15997 10839 16000
rect 10781 15991 10839 15997
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 11514 15960 11520 15972
rect 5684 15932 11520 15960
rect 5684 15920 5690 15932
rect 11514 15920 11520 15932
rect 11572 15920 11578 15972
rect 12406 15960 12434 16136
rect 17129 16133 17141 16167
rect 17175 16133 17187 16167
rect 18598 16164 18604 16176
rect 17129 16127 17187 16133
rect 17420 16136 18604 16164
rect 15654 16096 15660 16108
rect 15615 16068 15660 16096
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 17034 16096 17040 16108
rect 16995 16068 17040 16096
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 17310 16096 17316 16108
rect 17267 16068 17316 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17420 16105 17448 16136
rect 18598 16124 18604 16136
rect 18656 16124 18662 16176
rect 30282 16164 30288 16176
rect 18892 16136 30288 16164
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18121 16099 18179 16105
rect 18121 16096 18133 16099
rect 18012 16068 18133 16096
rect 18012 16056 18018 16068
rect 18121 16065 18133 16068
rect 18167 16065 18179 16099
rect 18121 16059 18179 16065
rect 14918 15988 14924 16040
rect 14976 16028 14982 16040
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 14976 16000 17877 16028
rect 14976 15988 14982 16000
rect 17865 15997 17877 16000
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 12406 15932 15608 15960
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 12710 15892 12716 15904
rect 10560 15864 12716 15892
rect 10560 15852 10566 15864
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 15470 15892 15476 15904
rect 15431 15864 15476 15892
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 15580 15892 15608 15932
rect 18892 15892 18920 16136
rect 30282 16124 30288 16136
rect 30340 16124 30346 16176
rect 21266 16096 21272 16108
rect 21227 16068 21272 16096
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 22261 16099 22319 16105
rect 22261 16096 22273 16099
rect 22112 16068 22273 16096
rect 22112 16028 22140 16068
rect 22261 16065 22273 16068
rect 22307 16065 22319 16099
rect 22261 16059 22319 16065
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16096 25191 16099
rect 25314 16096 25320 16108
rect 25179 16068 25320 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 25314 16056 25320 16068
rect 25372 16056 25378 16108
rect 27614 16096 27620 16108
rect 27575 16068 27620 16096
rect 27614 16056 27620 16068
rect 27672 16056 27678 16108
rect 27801 16099 27859 16105
rect 27801 16065 27813 16099
rect 27847 16065 27859 16099
rect 27801 16059 27859 16065
rect 28077 16099 28135 16105
rect 28077 16065 28089 16099
rect 28123 16065 28135 16099
rect 28077 16059 28135 16065
rect 28261 16099 28319 16105
rect 28261 16065 28273 16099
rect 28307 16096 28319 16099
rect 29181 16099 29239 16105
rect 29181 16096 29193 16099
rect 28307 16068 29193 16096
rect 28307 16065 28319 16068
rect 28261 16059 28319 16065
rect 29181 16065 29193 16068
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 21468 16000 22140 16028
rect 21468 15969 21496 16000
rect 23566 15988 23572 16040
rect 23624 16028 23630 16040
rect 24857 16031 24915 16037
rect 24857 16028 24869 16031
rect 23624 16000 24869 16028
rect 23624 15988 23630 16000
rect 24857 15997 24869 16000
rect 24903 15997 24915 16031
rect 24857 15991 24915 15997
rect 27430 15988 27436 16040
rect 27488 16028 27494 16040
rect 27816 16028 27844 16059
rect 27488 16000 27844 16028
rect 27488 15988 27494 16000
rect 21453 15963 21511 15969
rect 21453 15929 21465 15963
rect 21499 15929 21511 15963
rect 21453 15923 21511 15929
rect 27246 15920 27252 15972
rect 27304 15960 27310 15972
rect 28092 15960 28120 16059
rect 30098 16056 30104 16108
rect 30156 16096 30162 16108
rect 31113 16099 31171 16105
rect 31113 16096 31125 16099
rect 30156 16068 31125 16096
rect 30156 16056 30162 16068
rect 31113 16065 31125 16068
rect 31159 16065 31171 16099
rect 31113 16059 31171 16065
rect 31294 16056 31300 16108
rect 31352 16096 31358 16108
rect 36909 16099 36967 16105
rect 31352 16068 31445 16096
rect 31352 16056 31358 16068
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37734 16096 37740 16108
rect 36955 16068 37740 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 37734 16056 37740 16068
rect 37792 16056 37798 16108
rect 28905 16031 28963 16037
rect 28905 15997 28917 16031
rect 28951 15997 28963 16031
rect 28905 15991 28963 15997
rect 28997 16031 29055 16037
rect 28997 15997 29009 16031
rect 29043 15997 29055 16031
rect 28997 15991 29055 15997
rect 29089 16031 29147 16037
rect 29089 15997 29101 16031
rect 29135 16028 29147 16031
rect 30006 16028 30012 16040
rect 29135 16000 30012 16028
rect 29135 15997 29147 16000
rect 29089 15991 29147 15997
rect 27304 15932 28120 15960
rect 27304 15920 27310 15932
rect 28258 15920 28264 15972
rect 28316 15960 28322 15972
rect 28920 15960 28948 15991
rect 28316 15932 28948 15960
rect 29012 15960 29040 15991
rect 30006 15988 30012 16000
rect 30064 15988 30070 16040
rect 30193 16031 30251 16037
rect 30193 15997 30205 16031
rect 30239 16028 30251 16031
rect 30374 16028 30380 16040
rect 30239 16000 30380 16028
rect 30239 15997 30251 16000
rect 30193 15991 30251 15997
rect 30374 15988 30380 16000
rect 30432 15988 30438 16040
rect 30653 16031 30711 16037
rect 30653 15997 30665 16031
rect 30699 16028 30711 16031
rect 31312 16028 31340 16056
rect 30699 16000 31340 16028
rect 30699 15997 30711 16000
rect 30653 15991 30711 15997
rect 30561 15963 30619 15969
rect 29012 15932 30236 15960
rect 28316 15920 28322 15932
rect 30208 15904 30236 15932
rect 30561 15929 30573 15963
rect 30607 15960 30619 15963
rect 30926 15960 30932 15972
rect 30607 15932 30932 15960
rect 30607 15929 30619 15932
rect 30561 15923 30619 15929
rect 30926 15920 30932 15932
rect 30984 15920 30990 15972
rect 19242 15892 19248 15904
rect 15580 15864 18920 15892
rect 19203 15864 19248 15892
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 28718 15892 28724 15904
rect 28679 15864 28724 15892
rect 28718 15852 28724 15864
rect 28776 15852 28782 15904
rect 30190 15852 30196 15904
rect 30248 15892 30254 15904
rect 31113 15895 31171 15901
rect 31113 15892 31125 15895
rect 30248 15864 31125 15892
rect 30248 15852 30254 15864
rect 31113 15861 31125 15864
rect 31159 15861 31171 15895
rect 31113 15855 31171 15861
rect 36630 15852 36636 15904
rect 36688 15892 36694 15904
rect 36817 15895 36875 15901
rect 36817 15892 36829 15895
rect 36688 15864 36829 15892
rect 36688 15852 36694 15864
rect 36817 15861 36829 15864
rect 36863 15861 36875 15895
rect 37642 15892 37648 15904
rect 37603 15864 37648 15892
rect 36817 15855 36875 15861
rect 37642 15852 37648 15864
rect 37700 15852 37706 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 4706 15688 4712 15700
rect 4580 15660 4712 15688
rect 4580 15648 4586 15660
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 11422 15688 11428 15700
rect 9907 15660 11428 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 37458 15688 37464 15700
rect 11572 15660 37464 15688
rect 11572 15648 11578 15660
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 2222 15580 2228 15632
rect 2280 15620 2286 15632
rect 2280 15592 3464 15620
rect 2280 15580 2286 15592
rect 2866 15552 2872 15564
rect 2827 15524 2872 15552
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 3436 15561 3464 15592
rect 3421 15555 3479 15561
rect 3421 15521 3433 15555
rect 3467 15521 3479 15555
rect 3421 15515 3479 15521
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 10318 15552 10324 15564
rect 9723 15524 10324 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 11440 15552 11468 15648
rect 17954 15620 17960 15632
rect 17915 15592 17960 15620
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 23198 15620 23204 15632
rect 23159 15592 23204 15620
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 27982 15620 27988 15632
rect 26712 15592 27988 15620
rect 26712 15564 26740 15592
rect 27982 15580 27988 15592
rect 28040 15580 28046 15632
rect 30009 15623 30067 15629
rect 30009 15589 30021 15623
rect 30055 15589 30067 15623
rect 30558 15620 30564 15632
rect 30519 15592 30564 15620
rect 30009 15583 30067 15589
rect 14918 15552 14924 15564
rect 11440 15524 12664 15552
rect 14879 15524 14924 15552
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 9582 15484 9588 15496
rect 9543 15456 9588 15484
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 12636 15493 12664 15524
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 18230 15552 18236 15564
rect 17512 15524 18236 15552
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15484 12955 15487
rect 13722 15484 13728 15496
rect 12943 15456 13728 15484
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 3234 15416 3240 15428
rect 3195 15388 3240 15416
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 4249 15419 4307 15425
rect 4249 15385 4261 15419
rect 4295 15416 4307 15419
rect 4706 15416 4712 15428
rect 4295 15388 4712 15416
rect 4295 15385 4307 15388
rect 4249 15379 4307 15385
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 4264 15348 4292 15379
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 12452 15416 12480 15447
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 15188 15487 15246 15493
rect 15188 15453 15200 15487
rect 15234 15484 15246 15487
rect 15470 15484 15476 15496
rect 15234 15456 15476 15484
rect 15234 15453 15246 15456
rect 15188 15447 15246 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 17512 15493 17540 15524
rect 18230 15512 18236 15524
rect 18288 15512 18294 15564
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 22925 15555 22983 15561
rect 18748 15524 22094 15552
rect 18748 15512 18754 15524
rect 17313 15487 17371 15493
rect 17313 15484 17325 15487
rect 16264 15456 17325 15484
rect 16264 15444 16270 15456
rect 17313 15453 17325 15456
rect 17359 15453 17371 15487
rect 17313 15447 17371 15453
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 13538 15416 13544 15428
rect 12452 15388 13544 15416
rect 13538 15376 13544 15388
rect 13596 15376 13602 15428
rect 17034 15376 17040 15428
rect 17092 15416 17098 15428
rect 17604 15416 17632 15447
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 17736 15456 17781 15484
rect 17736 15444 17742 15456
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19300 15456 19533 15484
rect 19300 15444 19306 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 22066 15484 22094 15524
rect 22925 15521 22937 15555
rect 22971 15552 22983 15555
rect 23566 15552 23572 15564
rect 22971 15524 23572 15552
rect 22971 15521 22983 15524
rect 22925 15515 22983 15521
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 26694 15512 26700 15564
rect 26752 15552 26758 15564
rect 27430 15552 27436 15564
rect 26752 15524 26845 15552
rect 27391 15524 27436 15552
rect 26752 15512 26758 15524
rect 27430 15512 27436 15524
rect 27488 15512 27494 15564
rect 29086 15552 29092 15564
rect 29012 15524 29092 15552
rect 22833 15487 22891 15493
rect 22833 15484 22845 15487
rect 22066 15456 22845 15484
rect 19521 15447 19579 15453
rect 22833 15453 22845 15456
rect 22879 15453 22891 15487
rect 22833 15447 22891 15453
rect 27246 15444 27252 15496
rect 27304 15484 27310 15496
rect 29012 15493 29040 15524
rect 29086 15512 29092 15524
rect 29144 15512 29150 15564
rect 27341 15487 27399 15493
rect 27341 15484 27353 15487
rect 27304 15456 27353 15484
rect 27304 15444 27310 15456
rect 27341 15453 27353 15456
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15453 29055 15487
rect 28997 15447 29055 15453
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 30024 15484 30052 15583
rect 30558 15580 30564 15592
rect 30616 15580 30622 15632
rect 37642 15620 37648 15632
rect 36464 15592 37648 15620
rect 36464 15561 36492 15592
rect 37642 15580 37648 15592
rect 37700 15580 37706 15632
rect 36449 15555 36507 15561
rect 36449 15521 36461 15555
rect 36495 15521 36507 15555
rect 36630 15552 36636 15564
rect 36591 15524 36636 15552
rect 36449 15515 36507 15521
rect 36630 15512 36636 15524
rect 36688 15512 36694 15564
rect 38286 15552 38292 15564
rect 38247 15524 38292 15552
rect 38286 15512 38292 15524
rect 38344 15512 38350 15564
rect 29227 15456 30052 15484
rect 30190 15487 30248 15493
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 30190 15453 30202 15487
rect 30236 15484 30248 15487
rect 30374 15484 30380 15496
rect 30236 15456 30380 15484
rect 30236 15453 30248 15456
rect 30190 15447 30248 15453
rect 30374 15444 30380 15456
rect 30432 15444 30438 15496
rect 30650 15444 30656 15496
rect 30708 15484 30714 15496
rect 30708 15456 30753 15484
rect 30708 15444 30714 15456
rect 20070 15416 20076 15428
rect 17092 15388 20076 15416
rect 17092 15376 17098 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 26452 15419 26510 15425
rect 26452 15385 26464 15419
rect 26498 15416 26510 15419
rect 29089 15419 29147 15425
rect 29089 15416 29101 15419
rect 26498 15388 29101 15416
rect 26498 15385 26510 15388
rect 26452 15379 26510 15385
rect 29089 15385 29101 15388
rect 29135 15385 29147 15419
rect 29089 15379 29147 15385
rect 2372 15320 4292 15348
rect 2372 15308 2378 15320
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 9766 15348 9772 15360
rect 4856 15320 9772 15348
rect 4856 15308 4862 15320
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 12492 15320 13093 15348
rect 12492 15308 12498 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13081 15311 13139 15317
rect 16301 15351 16359 15357
rect 16301 15317 16313 15351
rect 16347 15348 16359 15351
rect 16482 15348 16488 15360
rect 16347 15320 16488 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 17586 15308 17592 15360
rect 17644 15348 17650 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 17644 15320 19625 15348
rect 17644 15308 17650 15320
rect 19613 15317 19625 15320
rect 19659 15348 19671 15351
rect 20162 15348 20168 15360
rect 19659 15320 20168 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 25317 15351 25375 15357
rect 25317 15317 25329 15351
rect 25363 15348 25375 15351
rect 25866 15348 25872 15360
rect 25363 15320 25872 15348
rect 25363 15317 25375 15320
rect 25317 15311 25375 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 27709 15351 27767 15357
rect 27709 15317 27721 15351
rect 27755 15348 27767 15351
rect 28258 15348 28264 15360
rect 27755 15320 28264 15348
rect 27755 15317 27767 15320
rect 27709 15311 27767 15317
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 30098 15308 30104 15360
rect 30156 15348 30162 15360
rect 30193 15351 30251 15357
rect 30193 15348 30205 15351
rect 30156 15320 30205 15348
rect 30156 15308 30162 15320
rect 30193 15317 30205 15320
rect 30239 15348 30251 15351
rect 30834 15348 30840 15360
rect 30239 15320 30840 15348
rect 30239 15317 30251 15320
rect 30193 15311 30251 15317
rect 30834 15308 30840 15320
rect 30892 15308 30898 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 12897 15147 12955 15153
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 13354 15144 13360 15156
rect 12943 15116 13360 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 19978 15144 19984 15156
rect 19208 15116 19984 15144
rect 19208 15104 19214 15116
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 20070 15104 20076 15156
rect 20128 15144 20134 15156
rect 21910 15144 21916 15156
rect 20128 15116 21916 15144
rect 20128 15104 20134 15116
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 23566 15144 23572 15156
rect 23527 15116 23572 15144
rect 23566 15104 23572 15116
rect 23624 15104 23630 15156
rect 26053 15147 26111 15153
rect 26053 15144 26065 15147
rect 24872 15116 26065 15144
rect 21266 15076 21272 15088
rect 19260 15048 21272 15076
rect 12434 15008 12440 15020
rect 12395 14980 12440 15008
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 12621 15014 12679 15017
rect 12621 15011 12848 15014
rect 12621 14977 12633 15011
rect 12667 15008 12848 15011
rect 13262 15008 13268 15020
rect 12667 14986 13268 15008
rect 12667 14977 12679 14986
rect 12820 14980 13268 14986
rect 12621 14971 12679 14977
rect 13262 14968 13268 14980
rect 13320 15008 13326 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 13320 14980 13369 15008
rect 13320 14968 13326 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13357 14971 13415 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 15008 14151 15011
rect 14182 15008 14188 15020
rect 14139 14980 14188 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 19260 15017 19288 15048
rect 21266 15036 21272 15048
rect 21324 15036 21330 15088
rect 24704 15079 24762 15085
rect 24704 15045 24716 15079
rect 24750 15076 24762 15079
rect 24872 15076 24900 15116
rect 26053 15113 26065 15116
rect 26099 15113 26111 15147
rect 30650 15144 30656 15156
rect 30611 15116 30656 15144
rect 26053 15107 26111 15113
rect 30650 15104 30656 15116
rect 30708 15104 30714 15156
rect 26694 15076 26700 15088
rect 24750 15048 24900 15076
rect 24964 15048 26700 15076
rect 24750 15045 24762 15048
rect 24704 15039 24762 15045
rect 24964 15020 24992 15048
rect 26694 15036 26700 15048
rect 26752 15036 26758 15088
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 14323 14980 19257 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 15008 19487 15011
rect 19475 14980 19932 15008
rect 19475 14977 19487 14980
rect 19429 14971 19487 14977
rect 1854 14940 1860 14952
rect 1815 14912 1860 14940
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2222 14940 2228 14952
rect 2087 14912 2228 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 12526 14940 12532 14952
rect 12584 14949 12590 14952
rect 2832 14912 2877 14940
rect 12495 14912 12532 14940
rect 2832 14900 2838 14912
rect 12526 14900 12532 14912
rect 12584 14903 12595 14949
rect 12584 14900 12590 14903
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 12768 14912 12813 14940
rect 12768 14900 12774 14912
rect 12728 14872 12756 14900
rect 14642 14872 14648 14884
rect 12728 14844 14648 14872
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 16114 14832 16120 14884
rect 16172 14872 16178 14884
rect 19904 14881 19932 14980
rect 19978 14968 19984 15020
rect 20036 15017 20042 15020
rect 20036 15011 20072 15017
rect 20060 15008 20072 15011
rect 21082 15008 21088 15020
rect 20060 14980 20668 15008
rect 21043 14980 21088 15008
rect 20060 14977 20072 14980
rect 20036 14971 20072 14977
rect 20036 14968 20042 14971
rect 20530 14940 20536 14952
rect 20491 14912 20536 14940
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 20640 14940 20668 14980
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 24946 15008 24952 15020
rect 24859 14980 24952 15008
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 15008 26203 15011
rect 27246 15008 27252 15020
rect 26191 14980 27252 15008
rect 26191 14977 26203 14980
rect 26145 14971 26203 14977
rect 21269 14943 21327 14949
rect 21269 14940 21281 14943
rect 20640 14912 21281 14940
rect 21269 14909 21281 14912
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 25976 14940 26004 14971
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 30282 15008 30288 15020
rect 30243 14980 30288 15008
rect 30282 14968 30288 14980
rect 30340 14968 30346 15020
rect 29086 14940 29092 14952
rect 25976 14912 29092 14940
rect 19889 14875 19947 14881
rect 16172 14844 19564 14872
rect 16172 14832 16178 14844
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 12860 14776 13461 14804
rect 12860 14764 12866 14776
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 14090 14804 14096 14816
rect 14051 14776 14096 14804
rect 13449 14767 13507 14773
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 19426 14804 19432 14816
rect 19387 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19536 14804 19564 14844
rect 19889 14841 19901 14875
rect 19935 14841 19947 14875
rect 19889 14835 19947 14841
rect 20441 14875 20499 14881
rect 20441 14841 20453 14875
rect 20487 14872 20499 14875
rect 22830 14872 22836 14884
rect 20487 14844 22836 14872
rect 20487 14841 20499 14844
rect 20441 14835 20499 14841
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 20990 14804 20996 14816
rect 19536 14776 20996 14804
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 25976 14804 26004 14912
rect 29086 14900 29092 14912
rect 29144 14900 29150 14952
rect 30190 14940 30196 14952
rect 30151 14912 30196 14940
rect 30190 14900 30196 14912
rect 30248 14900 30254 14952
rect 21324 14776 26004 14804
rect 21324 14764 21330 14776
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2685 14603 2743 14609
rect 2685 14569 2697 14603
rect 2731 14600 2743 14603
rect 3234 14600 3240 14612
rect 2731 14572 3240 14600
rect 2731 14569 2743 14572
rect 2685 14563 2743 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 16301 14603 16359 14609
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 16666 14600 16672 14612
rect 16347 14572 16672 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 18233 14603 18291 14609
rect 18233 14569 18245 14603
rect 18279 14600 18291 14603
rect 18414 14600 18420 14612
rect 18279 14572 18420 14600
rect 18279 14569 18291 14572
rect 18233 14563 18291 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19705 14603 19763 14609
rect 19705 14569 19717 14603
rect 19751 14600 19763 14603
rect 19978 14600 19984 14612
rect 19751 14572 19984 14600
rect 19751 14569 19763 14572
rect 19705 14563 19763 14569
rect 19978 14560 19984 14572
rect 20036 14600 20042 14612
rect 21082 14600 21088 14612
rect 20036 14572 21088 14600
rect 20036 14560 20042 14572
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 27246 14600 27252 14612
rect 27207 14572 27252 14600
rect 27246 14560 27252 14572
rect 27304 14560 27310 14612
rect 27614 14560 27620 14612
rect 27672 14600 27678 14612
rect 27801 14603 27859 14609
rect 27801 14600 27813 14603
rect 27672 14572 27813 14600
rect 27672 14560 27678 14572
rect 27801 14569 27813 14572
rect 27847 14569 27859 14603
rect 27801 14563 27859 14569
rect 28994 14560 29000 14612
rect 29052 14600 29058 14612
rect 30009 14603 30067 14609
rect 30009 14600 30021 14603
rect 29052 14572 30021 14600
rect 29052 14560 29058 14572
rect 30009 14569 30021 14572
rect 30055 14569 30067 14603
rect 30009 14563 30067 14569
rect 22370 14532 22376 14544
rect 22331 14504 22376 14532
rect 22370 14492 22376 14504
rect 22428 14492 22434 14544
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16224 14436 16865 14464
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 3050 14396 3056 14408
rect 2823 14368 3056 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 2884 14272 2912 14368
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10410 14396 10416 14408
rect 10367 14368 10416 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10410 14356 10416 14368
rect 10468 14356 10474 14408
rect 14918 14356 14924 14408
rect 14976 14396 14982 14408
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 14976 14368 15669 14396
rect 14976 14356 14982 14368
rect 15657 14365 15669 14368
rect 15703 14396 15715 14399
rect 16224 14396 16252 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 21085 14467 21143 14473
rect 21085 14433 21097 14467
rect 21131 14464 21143 14467
rect 22002 14464 22008 14476
rect 21131 14436 22008 14464
rect 21131 14433 21143 14436
rect 21085 14427 21143 14433
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 15703 14368 16252 14396
rect 15703 14365 15715 14368
rect 15657 14359 15715 14365
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16393 14399 16451 14405
rect 16393 14396 16405 14399
rect 16356 14368 16405 14396
rect 16356 14356 16362 14368
rect 16393 14365 16405 14368
rect 16439 14396 16451 14399
rect 16439 14368 19380 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 10226 14288 10232 14340
rect 10284 14328 10290 14340
rect 10566 14331 10624 14337
rect 10566 14328 10578 14331
rect 10284 14300 10578 14328
rect 10284 14288 10290 14300
rect 10566 14297 10578 14300
rect 10612 14297 10624 14331
rect 10566 14291 10624 14297
rect 14090 14288 14096 14340
rect 14148 14328 14154 14340
rect 15390 14331 15448 14337
rect 15390 14328 15402 14331
rect 14148 14300 15402 14328
rect 14148 14288 14154 14300
rect 15390 14297 15402 14300
rect 15436 14297 15448 14331
rect 15390 14291 15448 14297
rect 16206 14288 16212 14340
rect 16264 14328 16270 14340
rect 17098 14331 17156 14337
rect 17098 14328 17110 14331
rect 16264 14300 17110 14328
rect 16264 14288 16270 14300
rect 17098 14297 17110 14300
rect 17144 14297 17156 14331
rect 19352 14328 19380 14368
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 20818 14399 20876 14405
rect 20818 14396 20830 14399
rect 19484 14368 20830 14396
rect 19484 14356 19490 14368
rect 20818 14365 20830 14368
rect 20864 14365 20876 14399
rect 20818 14359 20876 14365
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 27430 14396 27436 14408
rect 22152 14368 22197 14396
rect 27391 14368 27436 14396
rect 22152 14356 22158 14368
rect 27430 14356 27436 14368
rect 27488 14356 27494 14408
rect 27890 14356 27896 14408
rect 27948 14396 27954 14408
rect 27948 14368 27993 14396
rect 27948 14356 27954 14368
rect 21818 14328 21824 14340
rect 19352 14300 21824 14328
rect 17098 14291 17156 14297
rect 21818 14288 21824 14300
rect 21876 14288 21882 14340
rect 22373 14331 22431 14337
rect 22373 14297 22385 14331
rect 22419 14328 22431 14331
rect 24854 14328 24860 14340
rect 22419 14300 24860 14328
rect 22419 14297 22431 14300
rect 22373 14291 22431 14297
rect 24854 14288 24860 14300
rect 24912 14328 24918 14340
rect 26510 14328 26516 14340
rect 24912 14300 26516 14328
rect 24912 14288 24918 14300
rect 26510 14288 26516 14300
rect 26568 14288 26574 14340
rect 29822 14288 29828 14340
rect 29880 14328 29886 14340
rect 29917 14331 29975 14337
rect 29917 14328 29929 14331
rect 29880 14300 29929 14328
rect 29880 14288 29886 14300
rect 29917 14297 29929 14300
rect 29963 14297 29975 14331
rect 29917 14291 29975 14297
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12710 14260 12716 14272
rect 11747 14232 12716 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 16114 14260 16120 14272
rect 16075 14232 16120 14260
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17586 14220 17592 14272
rect 17644 14260 17650 14272
rect 20070 14260 20076 14272
rect 17644 14232 20076 14260
rect 17644 14220 17650 14232
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 22186 14260 22192 14272
rect 22147 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 26326 14220 26332 14272
rect 26384 14260 26390 14272
rect 27433 14263 27491 14269
rect 27433 14260 27445 14263
rect 26384 14232 27445 14260
rect 26384 14220 26390 14232
rect 27433 14229 27445 14232
rect 27479 14260 27491 14263
rect 30098 14260 30104 14272
rect 27479 14232 30104 14260
rect 27479 14229 27491 14232
rect 27433 14223 27491 14229
rect 30098 14220 30104 14232
rect 30156 14220 30162 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 2222 14056 2228 14068
rect 2183 14028 2228 14056
rect 2222 14016 2228 14028
rect 2280 14016 2286 14068
rect 10226 14056 10232 14068
rect 10187 14028 10232 14056
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 12618 14056 12624 14068
rect 12579 14028 12624 14056
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 14182 14056 14188 14068
rect 14143 14028 14188 14056
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14642 14056 14648 14068
rect 14603 14028 14648 14056
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 16206 14056 16212 14068
rect 16167 14028 16212 14056
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 16298 14016 16304 14068
rect 16356 14016 16362 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19426 14056 19432 14068
rect 18739 14028 19432 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 19978 14056 19984 14068
rect 19843 14028 19984 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 20128 14028 20173 14056
rect 21284 14028 22109 14056
rect 20128 14016 20134 14028
rect 14553 13991 14611 13997
rect 14553 13957 14565 13991
rect 14599 13988 14611 13991
rect 15381 13991 15439 13997
rect 15381 13988 15393 13991
rect 14599 13960 15393 13988
rect 14599 13957 14611 13960
rect 14553 13951 14611 13957
rect 15381 13957 15393 13960
rect 15427 13957 15439 13991
rect 16316 13988 16344 14016
rect 19242 13988 19248 14000
rect 15381 13951 15439 13957
rect 15672 13960 16344 13988
rect 18984 13960 19248 13988
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 2314 13880 2320 13892
rect 2372 13920 2378 13932
rect 3142 13920 3148 13932
rect 2372 13892 3148 13920
rect 2372 13880 2378 13892
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 12710 13920 12716 13932
rect 12671 13892 12716 13920
rect 12710 13880 12716 13892
rect 12768 13920 12774 13932
rect 13538 13920 13544 13932
rect 12768 13892 13544 13920
rect 12768 13880 12774 13892
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14642 13880 14648 13932
rect 14700 13920 14706 13932
rect 14700 13892 15424 13920
rect 14700 13880 14706 13892
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15396 13861 15424 13892
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 15672 13929 15700 13960
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 15620 13892 15669 13920
rect 15620 13880 15626 13892
rect 15657 13889 15669 13892
rect 15703 13889 15715 13923
rect 16114 13920 16120 13932
rect 16075 13892 16120 13920
rect 15657 13883 15715 13889
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 16942 13920 16948 13932
rect 16347 13892 16948 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17218 13920 17224 13932
rect 17175 13892 17224 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 18984 13929 19012 13960
rect 19242 13948 19248 13960
rect 19300 13988 19306 14000
rect 21284 13997 21312 14028
rect 22097 14025 22109 14028
rect 22143 14025 22155 14059
rect 22097 14019 22155 14025
rect 25682 14016 25688 14068
rect 25740 14056 25746 14068
rect 25777 14059 25835 14065
rect 25777 14056 25789 14059
rect 25740 14028 25789 14056
rect 25740 14016 25746 14028
rect 25777 14025 25789 14028
rect 25823 14025 25835 14059
rect 27890 14056 27896 14068
rect 27851 14028 27896 14056
rect 25777 14019 25835 14025
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 19521 13991 19579 13997
rect 19521 13988 19533 13991
rect 19300 13960 19533 13988
rect 19300 13948 19306 13960
rect 19521 13957 19533 13960
rect 19567 13957 19579 13991
rect 19521 13951 19579 13957
rect 19889 13991 19947 13997
rect 19889 13957 19901 13991
rect 19935 13988 19947 13991
rect 21269 13991 21327 13997
rect 21269 13988 21281 13991
rect 19935 13960 21281 13988
rect 19935 13957 19947 13960
rect 19889 13951 19947 13957
rect 21269 13957 21281 13960
rect 21315 13957 21327 13991
rect 21269 13951 21327 13957
rect 22002 13948 22008 14000
rect 22060 13988 22066 14000
rect 24946 13988 24952 14000
rect 22060 13960 23520 13988
rect 22060 13948 22066 13960
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13889 19027 13923
rect 18969 13883 19027 13889
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13920 19119 13923
rect 19150 13920 19156 13932
rect 19107 13892 19156 13920
rect 19107 13889 19119 13892
rect 19061 13883 19119 13889
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13889 19763 13923
rect 19705 13883 19763 13889
rect 15381 13855 15439 13861
rect 14792 13824 14837 13852
rect 14792 13812 14798 13824
rect 15381 13821 15393 13855
rect 15427 13821 15439 13855
rect 15381 13815 15439 13821
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16540 13824 16865 13852
rect 16540 13812 16546 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 19720 13852 19748 13883
rect 22370 13880 22376 13932
rect 22428 13920 22434 13932
rect 23492 13929 23520 13960
rect 24412 13960 24952 13988
rect 24412 13929 24440 13960
rect 24946 13948 24952 13960
rect 25004 13948 25010 14000
rect 23210 13923 23268 13929
rect 23210 13920 23222 13923
rect 22428 13892 23222 13920
rect 22428 13880 22434 13892
rect 23210 13889 23222 13892
rect 23256 13889 23268 13923
rect 23210 13883 23268 13889
rect 23477 13923 23535 13929
rect 23477 13889 23489 13923
rect 23523 13920 23535 13923
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 23523 13892 24409 13920
rect 23523 13889 23535 13892
rect 23477 13883 23535 13889
rect 24397 13889 24409 13892
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 24664 13923 24722 13929
rect 24664 13889 24676 13923
rect 24710 13920 24722 13923
rect 25130 13920 25136 13932
rect 24710 13892 25136 13920
rect 24710 13889 24722 13892
rect 24664 13883 24722 13889
rect 25130 13880 25136 13892
rect 25188 13880 25194 13932
rect 27982 13880 27988 13932
rect 28040 13920 28046 13932
rect 28261 13923 28319 13929
rect 28261 13920 28273 13923
rect 28040 13892 28273 13920
rect 28040 13880 28046 13892
rect 28261 13889 28273 13892
rect 28307 13889 28319 13923
rect 29178 13920 29184 13932
rect 29139 13892 29184 13920
rect 28261 13883 28319 13889
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13920 29423 13923
rect 29822 13920 29828 13932
rect 29411 13892 29828 13920
rect 29411 13889 29423 13892
rect 29365 13883 29423 13889
rect 29822 13880 29828 13892
rect 29880 13880 29886 13932
rect 30098 13920 30104 13932
rect 30059 13892 30104 13920
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 16853 13815 16911 13821
rect 18892 13824 19748 13852
rect 21453 13855 21511 13861
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 12618 13784 12624 13796
rect 9180 13756 12624 13784
rect 9180 13744 9186 13756
rect 12618 13744 12624 13756
rect 12676 13744 12682 13796
rect 15565 13787 15623 13793
rect 15565 13753 15577 13787
rect 15611 13784 15623 13787
rect 16666 13784 16672 13796
rect 15611 13756 16672 13784
rect 15611 13753 15623 13756
rect 15565 13747 15623 13753
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 18892 13725 18920 13824
rect 21453 13821 21465 13855
rect 21499 13852 21511 13855
rect 21499 13824 22094 13852
rect 21499 13821 21511 13824
rect 21453 13815 21511 13821
rect 18877 13719 18935 13725
rect 18877 13716 18889 13719
rect 18472 13688 18889 13716
rect 18472 13676 18478 13688
rect 18877 13685 18889 13688
rect 18923 13685 18935 13719
rect 22066 13716 22094 13824
rect 28074 13812 28080 13864
rect 28132 13852 28138 13864
rect 28353 13855 28411 13861
rect 28353 13852 28365 13855
rect 28132 13824 28365 13852
rect 28132 13812 28138 13824
rect 28353 13821 28365 13824
rect 28399 13852 28411 13855
rect 28718 13852 28724 13864
rect 28399 13824 28724 13852
rect 28399 13821 28411 13824
rect 28353 13815 28411 13821
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 28997 13855 29055 13861
rect 28997 13821 29009 13855
rect 29043 13852 29055 13855
rect 29914 13852 29920 13864
rect 29043 13824 29920 13852
rect 29043 13821 29055 13824
rect 28997 13815 29055 13821
rect 29914 13812 29920 13824
rect 29972 13812 29978 13864
rect 22738 13716 22744 13728
rect 22066 13688 22744 13716
rect 18877 13679 18935 13685
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 10042 13512 10048 13524
rect 9999 13484 10048 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10318 13472 10324 13524
rect 10376 13512 10382 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 10376 13484 12633 13512
rect 10376 13472 10382 13484
rect 12621 13481 12633 13484
rect 12667 13512 12679 13515
rect 13262 13512 13268 13524
rect 12667 13484 13268 13512
rect 12667 13481 12679 13484
rect 12621 13475 12679 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13357 13515 13415 13521
rect 13357 13481 13369 13515
rect 13403 13512 13415 13515
rect 14734 13512 14740 13524
rect 13403 13484 14740 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17865 13515 17923 13521
rect 17865 13481 17877 13515
rect 17911 13512 17923 13515
rect 18506 13512 18512 13524
rect 17911 13484 18512 13512
rect 17911 13481 17923 13484
rect 17865 13475 17923 13481
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 21910 13512 21916 13524
rect 21871 13484 21916 13512
rect 21910 13472 21916 13484
rect 21968 13512 21974 13524
rect 21968 13484 22094 13512
rect 21968 13472 21974 13484
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 12802 13444 12808 13456
rect 12584 13416 12808 13444
rect 12584 13404 12590 13416
rect 12802 13404 12808 13416
rect 12860 13404 12866 13456
rect 16666 13404 16672 13456
rect 16724 13444 16730 13456
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 16724 13416 17049 13444
rect 16724 13404 16730 13416
rect 17037 13413 17049 13416
rect 17083 13413 17095 13447
rect 17037 13407 17095 13413
rect 10410 13376 10416 13388
rect 10371 13348 10416 13376
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 17954 13376 17960 13388
rect 16899 13348 17960 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 22066 13376 22094 13484
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22244 13484 22845 13512
rect 22244 13472 22250 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 23750 13512 23756 13524
rect 23711 13484 23756 13512
rect 22833 13475 22891 13481
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 25130 13512 25136 13524
rect 25091 13484 25136 13512
rect 25130 13472 25136 13484
rect 25188 13472 25194 13524
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 26697 13515 26755 13521
rect 25740 13484 26280 13512
rect 25740 13472 25746 13484
rect 26145 13447 26203 13453
rect 26145 13413 26157 13447
rect 26191 13413 26203 13447
rect 26145 13407 26203 13413
rect 22066 13348 22968 13376
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 12250 13308 12256 13320
rect 11296 13280 12256 13308
rect 11296 13268 11302 13280
rect 12250 13268 12256 13280
rect 12308 13308 12314 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 12308 13280 13185 13308
rect 12308 13268 12314 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 13173 13271 13231 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17552 13280 17601 13308
rect 17552 13268 17558 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 21818 13268 21824 13320
rect 21876 13308 21882 13320
rect 22097 13311 22155 13317
rect 22097 13308 22109 13311
rect 21876 13280 22109 13308
rect 21876 13268 21882 13280
rect 22097 13277 22109 13280
rect 22143 13277 22155 13311
rect 22097 13271 22155 13277
rect 22281 13311 22339 13317
rect 22281 13277 22293 13311
rect 22327 13277 22339 13311
rect 22738 13308 22744 13320
rect 22699 13280 22744 13308
rect 22281 13271 22339 13277
rect 9490 13200 9496 13252
rect 9548 13240 9554 13252
rect 9585 13243 9643 13249
rect 9585 13240 9597 13243
rect 9548 13212 9597 13240
rect 9548 13200 9554 13212
rect 9585 13209 9597 13212
rect 9631 13209 9643 13243
rect 9585 13203 9643 13209
rect 9769 13243 9827 13249
rect 9769 13209 9781 13243
rect 9815 13240 9827 13243
rect 10410 13240 10416 13252
rect 9815 13212 10416 13240
rect 9815 13209 9827 13212
rect 9769 13203 9827 13209
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 10686 13249 10692 13252
rect 10680 13240 10692 13249
rect 10647 13212 10692 13240
rect 10680 13203 10692 13212
rect 10686 13200 10692 13203
rect 10744 13200 10750 13252
rect 12529 13243 12587 13249
rect 12529 13240 12541 13243
rect 12406 13212 12541 13240
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 12406 13172 12434 13212
rect 12529 13209 12541 13212
rect 12575 13240 12587 13243
rect 14182 13240 14188 13252
rect 12575 13212 14188 13240
rect 12575 13209 12587 13212
rect 12529 13203 12587 13209
rect 14182 13200 14188 13212
rect 14240 13200 14246 13252
rect 17770 13200 17776 13252
rect 17828 13240 17834 13252
rect 22296 13240 22324 13271
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 22940 13317 22968 13348
rect 22925 13311 22983 13317
rect 22925 13277 22937 13311
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 24854 13268 24860 13320
rect 24912 13308 24918 13320
rect 24949 13311 25007 13317
rect 24949 13308 24961 13311
rect 24912 13280 24961 13308
rect 24912 13268 24918 13280
rect 24949 13277 24961 13280
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13308 25191 13311
rect 26160 13308 26188 13407
rect 25179 13280 26188 13308
rect 26252 13317 26280 13484
rect 26697 13481 26709 13515
rect 26743 13512 26755 13515
rect 27522 13512 27528 13524
rect 26743 13484 27528 13512
rect 26743 13481 26755 13484
rect 26697 13475 26755 13481
rect 27522 13472 27528 13484
rect 27580 13472 27586 13524
rect 26252 13311 26328 13317
rect 26252 13280 26282 13311
rect 25179 13277 25191 13280
rect 25133 13271 25191 13277
rect 26270 13277 26282 13280
rect 26316 13277 26328 13311
rect 26270 13271 26328 13277
rect 26786 13268 26792 13320
rect 26844 13308 26850 13320
rect 27798 13308 27804 13320
rect 26844 13280 26889 13308
rect 27759 13280 27804 13308
rect 26844 13268 26850 13280
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 28074 13308 28080 13320
rect 28035 13280 28080 13308
rect 28074 13268 28080 13280
rect 28132 13268 28138 13320
rect 37829 13311 37887 13317
rect 37829 13277 37841 13311
rect 37875 13308 37887 13311
rect 38286 13308 38292 13320
rect 37875 13280 38292 13308
rect 37875 13277 37887 13280
rect 37829 13271 37887 13277
rect 38286 13268 38292 13280
rect 38344 13268 38350 13320
rect 23845 13243 23903 13249
rect 23845 13240 23857 13243
rect 17828 13212 17873 13240
rect 22296 13212 23857 13240
rect 17828 13200 17834 13212
rect 23845 13209 23857 13212
rect 23891 13240 23903 13243
rect 29914 13240 29920 13252
rect 23891 13212 29920 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 29914 13200 29920 13212
rect 29972 13200 29978 13252
rect 26326 13172 26332 13184
rect 11839 13144 12434 13172
rect 26287 13144 26332 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 26326 13132 26332 13144
rect 26384 13132 26390 13184
rect 27614 13172 27620 13184
rect 27575 13144 27620 13172
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 27982 13172 27988 13184
rect 27943 13144 27988 13172
rect 27982 13132 27988 13144
rect 28040 13132 28046 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 10318 12968 10324 12980
rect 10279 12940 10324 12968
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 14182 12928 14188 12980
rect 14240 12968 14246 12980
rect 15381 12971 15439 12977
rect 15381 12968 15393 12971
rect 14240 12940 15393 12968
rect 14240 12928 14246 12940
rect 15381 12937 15393 12940
rect 15427 12937 15439 12971
rect 15381 12931 15439 12937
rect 17313 12971 17371 12977
rect 17313 12937 17325 12971
rect 17359 12968 17371 12971
rect 17494 12968 17500 12980
rect 17359 12940 17500 12968
rect 17359 12937 17371 12940
rect 17313 12931 17371 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 17954 12968 17960 12980
rect 17915 12940 17960 12968
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 19242 12928 19248 12980
rect 19300 12968 19306 12980
rect 20162 12968 20168 12980
rect 19300 12940 20168 12968
rect 19300 12928 19306 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 26513 12971 26571 12977
rect 26513 12937 26525 12971
rect 26559 12968 26571 12971
rect 26786 12968 26792 12980
rect 26559 12940 26792 12968
rect 26559 12937 26571 12940
rect 26513 12931 26571 12937
rect 26786 12928 26792 12940
rect 26844 12928 26850 12980
rect 27798 12968 27804 12980
rect 27759 12940 27804 12968
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 10686 12900 10692 12912
rect 10647 12872 10692 12900
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 14274 12860 14280 12912
rect 14332 12900 14338 12912
rect 14642 12900 14648 12912
rect 14332 12872 14648 12900
rect 14332 12860 14338 12872
rect 14642 12860 14648 12872
rect 14700 12900 14706 12912
rect 14737 12903 14795 12909
rect 14737 12900 14749 12903
rect 14700 12872 14749 12900
rect 14700 12860 14706 12872
rect 14737 12869 14749 12872
rect 14783 12869 14795 12903
rect 15565 12903 15623 12909
rect 15565 12900 15577 12903
rect 14737 12863 14795 12869
rect 14844 12872 15577 12900
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 2314 12832 2320 12844
rect 2271 12804 2320 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 9122 12832 9128 12844
rect 9083 12804 9128 12832
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 10226 12832 10232 12844
rect 10187 12804 10232 12832
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10468 12804 10609 12832
rect 10468 12792 10474 12804
rect 10597 12801 10609 12804
rect 10643 12832 10655 12835
rect 13265 12835 13323 12841
rect 10643 12804 13216 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 11238 12764 11244 12776
rect 9263 12736 11244 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12768 12736 13001 12764
rect 12768 12724 12774 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 13188 12764 13216 12804
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 13998 12832 14004 12844
rect 13311 12804 14004 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13998 12792 14004 12804
rect 14056 12832 14062 12844
rect 14844 12832 14872 12872
rect 15565 12869 15577 12872
rect 15611 12869 15623 12903
rect 16482 12900 16488 12912
rect 15565 12863 15623 12869
rect 16040 12872 16488 12900
rect 15286 12832 15292 12844
rect 14056 12804 14872 12832
rect 15247 12804 15292 12832
rect 14056 12792 14062 12804
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15654 12792 15660 12844
rect 15712 12832 15718 12844
rect 16040 12841 16068 12872
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 17586 12900 17592 12912
rect 17144 12872 17592 12900
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15712 12804 16037 12832
rect 15712 12792 15718 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12832 16267 12835
rect 17144 12832 17172 12872
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 17770 12860 17776 12912
rect 17828 12900 17834 12912
rect 19521 12903 19579 12909
rect 17828 12872 18552 12900
rect 17828 12860 17834 12872
rect 16255 12804 17172 12832
rect 17221 12835 17279 12841
rect 16255 12801 16267 12804
rect 16209 12795 16267 12801
rect 17221 12801 17233 12835
rect 17267 12801 17279 12835
rect 17402 12832 17408 12844
rect 17363 12804 17408 12832
rect 17221 12795 17279 12801
rect 16114 12764 16120 12776
rect 13188 12736 16120 12764
rect 12989 12727 13047 12733
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 9950 12696 9956 12708
rect 4120 12668 9956 12696
rect 4120 12656 4126 12668
rect 9950 12656 9956 12668
rect 10008 12656 10014 12708
rect 13004 12696 13032 12727
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 17236 12764 17264 12795
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 18138 12832 18144 12844
rect 18099 12804 18144 12832
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18414 12832 18420 12844
rect 18288 12804 18333 12832
rect 18375 12804 18420 12832
rect 18288 12792 18294 12804
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18524 12841 18552 12872
rect 19521 12869 19533 12903
rect 19567 12900 19579 12903
rect 29178 12900 29184 12912
rect 19567 12872 20300 12900
rect 19567 12869 19579 12872
rect 19521 12863 19579 12869
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12801 18567 12835
rect 19242 12832 19248 12844
rect 19203 12804 19248 12832
rect 18509 12795 18567 12801
rect 16224 12736 17264 12764
rect 16224 12708 16252 12736
rect 13446 12696 13452 12708
rect 13004 12668 13452 12696
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 14550 12696 14556 12708
rect 14511 12668 14556 12696
rect 14550 12656 14556 12668
rect 14608 12696 14614 12708
rect 15286 12696 15292 12708
rect 14608 12668 15292 12696
rect 14608 12656 14614 12668
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 15565 12699 15623 12705
rect 15565 12665 15577 12699
rect 15611 12696 15623 12699
rect 16206 12696 16212 12708
rect 15611 12668 16212 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 18524 12696 18552 12795
rect 19242 12792 19248 12804
rect 19300 12792 19306 12844
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 20162 12832 20168 12844
rect 19484 12804 20168 12832
rect 19484 12792 19490 12804
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20272 12841 20300 12872
rect 22066 12872 29184 12900
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12801 20315 12835
rect 20257 12795 20315 12801
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 19392 12736 19533 12764
rect 19392 12724 19398 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 22066 12696 22094 12872
rect 29178 12860 29184 12872
rect 29236 12860 29242 12912
rect 25133 12835 25191 12841
rect 25133 12801 25145 12835
rect 25179 12801 25191 12835
rect 25682 12832 25688 12844
rect 25133 12795 25191 12801
rect 25240 12804 25688 12832
rect 18524 12668 22094 12696
rect 25148 12696 25176 12795
rect 25240 12773 25268 12804
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 26145 12835 26203 12841
rect 26145 12801 26157 12835
rect 26191 12832 26203 12835
rect 27614 12832 27620 12844
rect 26191 12804 27620 12832
rect 26191 12801 26203 12804
rect 26145 12795 26203 12801
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 37461 12835 37519 12841
rect 37461 12801 37473 12835
rect 37507 12832 37519 12835
rect 37918 12832 37924 12844
rect 37507 12804 37924 12832
rect 37507 12801 37519 12804
rect 37461 12795 37519 12801
rect 37918 12792 37924 12804
rect 37976 12792 37982 12844
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12733 25283 12767
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25225 12727 25283 12733
rect 25516 12736 26065 12764
rect 25516 12705 25544 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 27154 12724 27160 12776
rect 27212 12764 27218 12776
rect 27341 12767 27399 12773
rect 27341 12764 27353 12767
rect 27212 12736 27353 12764
rect 27212 12724 27218 12736
rect 27341 12733 27353 12736
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 27430 12724 27436 12776
rect 27488 12764 27494 12776
rect 28721 12767 28779 12773
rect 28721 12764 28733 12767
rect 27488 12736 28733 12764
rect 27488 12724 27494 12736
rect 25501 12699 25559 12705
rect 25148 12668 25268 12696
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 1820 12600 2145 12628
rect 1820 12588 1826 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 10502 12628 10508 12640
rect 10463 12600 10508 12628
rect 2133 12591 2191 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 12710 12628 12716 12640
rect 12671 12600 12716 12628
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13173 12631 13231 12637
rect 13173 12597 13185 12631
rect 13219 12628 13231 12631
rect 13262 12628 13268 12640
rect 13219 12600 13268 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 15746 12588 15752 12640
rect 15804 12628 15810 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15804 12600 16129 12628
rect 15804 12588 15810 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 19150 12628 19156 12640
rect 17184 12600 19156 12628
rect 17184 12588 17190 12600
rect 19150 12588 19156 12600
rect 19208 12628 19214 12640
rect 19337 12631 19395 12637
rect 19337 12628 19349 12631
rect 19208 12600 19349 12628
rect 19208 12588 19214 12600
rect 19337 12597 19349 12600
rect 19383 12597 19395 12631
rect 19978 12628 19984 12640
rect 19939 12600 19984 12628
rect 19337 12591 19395 12597
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 25240 12628 25268 12668
rect 25501 12665 25513 12699
rect 25547 12665 25559 12699
rect 25501 12659 25559 12665
rect 27172 12628 27200 12724
rect 27724 12705 27752 12736
rect 28721 12733 28733 12736
rect 28767 12733 28779 12767
rect 28721 12727 28779 12733
rect 27709 12699 27767 12705
rect 27709 12665 27721 12699
rect 27755 12665 27767 12699
rect 28353 12699 28411 12705
rect 28353 12696 28365 12699
rect 27709 12659 27767 12665
rect 27816 12668 28365 12696
rect 27816 12628 27844 12668
rect 28353 12665 28365 12668
rect 28399 12665 28411 12699
rect 28353 12659 28411 12665
rect 25240 12600 27844 12628
rect 28074 12588 28080 12640
rect 28132 12628 28138 12640
rect 28261 12631 28319 12637
rect 28261 12628 28273 12631
rect 28132 12600 28273 12628
rect 28132 12588 28138 12600
rect 28261 12597 28273 12600
rect 28307 12597 28319 12631
rect 28261 12591 28319 12597
rect 37553 12631 37611 12637
rect 37553 12597 37565 12631
rect 37599 12628 37611 12631
rect 38102 12628 38108 12640
rect 37599 12600 38108 12628
rect 37599 12597 37611 12600
rect 37553 12591 37611 12597
rect 38102 12588 38108 12600
rect 38160 12588 38166 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 10560 12396 10609 12424
rect 10560 12384 10566 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13354 12424 13360 12436
rect 13035 12396 13360 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 13504 12396 14473 12424
rect 13504 12384 13510 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 14461 12387 14519 12393
rect 16577 12427 16635 12433
rect 16577 12393 16589 12427
rect 16623 12424 16635 12427
rect 17310 12424 17316 12436
rect 16623 12396 17316 12424
rect 16623 12393 16635 12396
rect 16577 12387 16635 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18233 12427 18291 12433
rect 18233 12393 18245 12427
rect 18279 12424 18291 12427
rect 18414 12424 18420 12436
rect 18279 12396 18420 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20441 12427 20499 12433
rect 20441 12393 20453 12427
rect 20487 12424 20499 12427
rect 20530 12424 20536 12436
rect 20487 12396 20536 12424
rect 20487 12393 20499 12396
rect 20441 12387 20499 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 21910 12424 21916 12436
rect 21871 12396 21916 12424
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 22094 12424 22100 12436
rect 22055 12396 22100 12424
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 27982 12384 27988 12436
rect 28040 12424 28046 12436
rect 28077 12427 28135 12433
rect 28077 12424 28089 12427
rect 28040 12396 28089 12424
rect 28040 12384 28046 12396
rect 28077 12393 28089 12396
rect 28123 12393 28135 12427
rect 28077 12387 28135 12393
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14553 12359 14611 12365
rect 14553 12356 14565 12359
rect 14240 12328 14565 12356
rect 14240 12316 14246 12328
rect 14553 12325 14565 12328
rect 14599 12325 14611 12359
rect 14553 12319 14611 12325
rect 15013 12359 15071 12365
rect 15013 12325 15025 12359
rect 15059 12356 15071 12359
rect 15562 12356 15568 12368
rect 15059 12328 15568 12356
rect 15059 12325 15071 12328
rect 15013 12319 15071 12325
rect 15562 12316 15568 12328
rect 15620 12356 15626 12368
rect 17402 12356 17408 12368
rect 15620 12328 17408 12356
rect 15620 12316 15626 12328
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 18138 12316 18144 12368
rect 18196 12356 18202 12368
rect 18785 12359 18843 12365
rect 18785 12356 18797 12359
rect 18196 12328 18797 12356
rect 18196 12316 18202 12328
rect 18785 12325 18797 12328
rect 18831 12325 18843 12359
rect 18785 12319 18843 12325
rect 21177 12359 21235 12365
rect 21177 12325 21189 12359
rect 21223 12325 21235 12359
rect 21177 12319 21235 12325
rect 1762 12288 1768 12300
rect 1723 12260 1768 12288
rect 1762 12248 1768 12260
rect 1820 12248 1826 12300
rect 2774 12288 2780 12300
rect 2735 12260 2780 12288
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 10226 12248 10232 12300
rect 10284 12288 10290 12300
rect 11609 12291 11667 12297
rect 11609 12288 11621 12291
rect 10284 12260 11621 12288
rect 10284 12248 10290 12260
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 10318 12180 10324 12232
rect 10376 12220 10382 12232
rect 10612 12229 10640 12260
rect 11609 12257 11621 12260
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12342 12288 12348 12300
rect 11747 12260 12348 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12526 12288 12532 12300
rect 12487 12260 12532 12288
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 12894 12288 12900 12300
rect 12667 12260 12900 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 15654 12288 15660 12300
rect 14292 12260 15660 12288
rect 10413 12223 10471 12229
rect 10413 12220 10425 12223
rect 10376 12192 10425 12220
rect 10376 12180 10382 12192
rect 10413 12189 10425 12192
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 11848 12192 11893 12220
rect 11848 12180 11854 12192
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 14292 12229 14320 12260
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 15804 12260 16313 12288
rect 15804 12248 15810 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 17420 12288 17448 12316
rect 18800 12288 18828 12319
rect 21192 12288 21220 12319
rect 37182 12288 37188 12300
rect 17420 12260 18736 12288
rect 18800 12260 19932 12288
rect 16301 12251 16359 12257
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 12768 12192 12817 12220
rect 12768 12180 12774 12192
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14642 12220 14648 12232
rect 14603 12192 14648 12220
rect 14277 12183 14335 12189
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 14734 12180 14740 12232
rect 14792 12220 14798 12232
rect 16114 12220 16120 12232
rect 14792 12192 14837 12220
rect 16075 12192 16120 12220
rect 14792 12180 14798 12192
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 16393 12223 16451 12229
rect 16264 12192 16309 12220
rect 16264 12180 16270 12192
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 16439 12192 17049 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 17037 12189 17049 12192
rect 17083 12189 17095 12223
rect 17218 12220 17224 12232
rect 17179 12192 17224 12220
rect 17037 12183 17095 12189
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 17586 12220 17592 12232
rect 17451 12192 17592 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 12069 12155 12127 12161
rect 12069 12121 12081 12155
rect 12115 12152 12127 12155
rect 12526 12152 12532 12164
rect 12115 12124 12532 12152
rect 12115 12121 12127 12124
rect 12069 12115 12127 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 11974 12084 11980 12096
rect 11887 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12084 12038 12096
rect 12618 12084 12624 12096
rect 12032 12056 12624 12084
rect 12032 12044 12038 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 16206 12044 16212 12096
rect 16264 12084 16270 12096
rect 18064 12084 18092 12183
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 18414 12220 18420 12232
rect 18288 12192 18420 12220
rect 18288 12180 18294 12192
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 18708 12229 18736 12260
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12189 18751 12223
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18693 12183 18751 12189
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19904 12229 19932 12260
rect 20180 12260 21220 12288
rect 37143 12260 37188 12288
rect 20180 12229 20208 12260
rect 37182 12248 37188 12260
rect 37240 12248 37246 12300
rect 38102 12288 38108 12300
rect 38063 12260 38108 12288
rect 38102 12248 38108 12260
rect 38160 12248 38166 12300
rect 38286 12288 38292 12300
rect 38247 12260 38292 12288
rect 38286 12248 38292 12260
rect 38344 12248 38350 12300
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20898 12220 20904 12232
rect 20312 12192 20357 12220
rect 20859 12192 20904 12220
rect 20312 12180 20318 12192
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 21508 12192 21741 12220
rect 21508 12180 21514 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 21876 12192 21921 12220
rect 21876 12180 21882 12192
rect 27798 12180 27804 12232
rect 27856 12220 27862 12232
rect 27893 12223 27951 12229
rect 27893 12220 27905 12223
rect 27856 12192 27905 12220
rect 27856 12180 27862 12192
rect 27893 12189 27905 12192
rect 27939 12189 27951 12223
rect 28074 12220 28080 12232
rect 28035 12192 28080 12220
rect 27893 12183 27951 12189
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 19426 12112 19432 12164
rect 19484 12152 19490 12164
rect 20070 12152 20076 12164
rect 19484 12124 20076 12152
rect 19484 12112 19490 12124
rect 20070 12112 20076 12124
rect 20128 12152 20134 12164
rect 21177 12155 21235 12161
rect 21177 12152 21189 12155
rect 20128 12124 21189 12152
rect 20128 12112 20134 12124
rect 21177 12121 21189 12124
rect 21223 12121 21235 12155
rect 21177 12115 21235 12121
rect 16264 12056 18092 12084
rect 16264 12044 16270 12056
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 20993 12087 21051 12093
rect 20993 12084 21005 12087
rect 19392 12056 21005 12084
rect 19392 12044 19398 12056
rect 20993 12053 21005 12056
rect 21039 12053 21051 12087
rect 20993 12047 21051 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 11977 11883 12035 11889
rect 11977 11849 11989 11883
rect 12023 11880 12035 11883
rect 12894 11880 12900 11892
rect 12023 11852 12900 11880
rect 12023 11849 12035 11852
rect 11977 11843 12035 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 16172 11852 16313 11880
rect 16172 11840 16178 11852
rect 16301 11849 16313 11852
rect 16347 11849 16359 11883
rect 16301 11843 16359 11849
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17368 11852 21496 11880
rect 17368 11840 17374 11852
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 14921 11815 14979 11821
rect 12584 11784 13216 11812
rect 12584 11772 12590 11784
rect 1578 11704 1584 11756
rect 1636 11744 1642 11756
rect 1857 11747 1915 11753
rect 1857 11744 1869 11747
rect 1636 11716 1869 11744
rect 1636 11704 1642 11716
rect 1857 11713 1869 11716
rect 1903 11713 1915 11747
rect 1857 11707 1915 11713
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9824 11716 9965 11744
rect 9824 11704 9830 11716
rect 9953 11713 9965 11716
rect 9999 11744 10011 11747
rect 10502 11744 10508 11756
rect 9999 11716 10508 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 11974 11744 11980 11756
rect 11839 11716 11980 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11744 12127 11747
rect 12805 11747 12863 11753
rect 12115 11716 12756 11744
rect 12115 11713 12127 11716
rect 12069 11707 12127 11713
rect 12728 11685 12756 11716
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 12851 11716 13124 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 12713 11679 12771 11685
rect 12713 11645 12725 11679
rect 12759 11676 12771 11679
rect 12759 11648 13032 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 11790 11608 11796 11620
rect 11751 11580 11796 11608
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 10045 11543 10103 11549
rect 10045 11509 10057 11543
rect 10091 11540 10103 11543
rect 11606 11540 11612 11552
rect 10091 11512 11612 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 12529 11543 12587 11549
rect 12529 11509 12541 11543
rect 12575 11540 12587 11543
rect 12710 11540 12716 11552
rect 12575 11512 12716 11540
rect 12575 11509 12587 11512
rect 12529 11503 12587 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 13004 11540 13032 11648
rect 13096 11608 13124 11716
rect 13188 11685 13216 11784
rect 14921 11781 14933 11815
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 15105 11815 15163 11821
rect 15105 11781 15117 11815
rect 15151 11812 15163 11815
rect 15746 11812 15752 11824
rect 15151 11784 15752 11812
rect 15151 11781 15163 11784
rect 15105 11775 15163 11781
rect 13998 11744 14004 11756
rect 13959 11716 14004 11744
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11744 14335 11747
rect 14642 11744 14648 11756
rect 14323 11716 14648 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 14737 11679 14795 11685
rect 14737 11676 14749 11679
rect 13219 11648 14749 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 14737 11645 14749 11648
rect 14783 11645 14795 11679
rect 14737 11639 14795 11645
rect 13817 11611 13875 11617
rect 13817 11608 13829 11611
rect 13096 11580 13829 11608
rect 13817 11577 13829 11580
rect 13863 11608 13875 11611
rect 14458 11608 14464 11620
rect 13863 11580 14464 11608
rect 13863 11577 13875 11580
rect 13817 11571 13875 11577
rect 14458 11568 14464 11580
rect 14516 11608 14522 11620
rect 14936 11608 14964 11775
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 18874 11812 18880 11824
rect 15856 11784 18880 11812
rect 15856 11756 15884 11784
rect 18874 11772 18880 11784
rect 18932 11812 18938 11824
rect 18932 11784 19748 11812
rect 18932 11772 18938 11784
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 15620 11716 15669 11744
rect 15620 11704 15626 11716
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 15838 11744 15844 11756
rect 15751 11716 15844 11744
rect 15657 11707 15715 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16206 11744 16212 11756
rect 16071 11716 16212 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 15948 11676 15976 11707
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11742 18107 11747
rect 19334 11744 19340 11756
rect 18136 11742 19196 11744
rect 18095 11716 19196 11742
rect 19247 11716 19340 11744
rect 18095 11714 18164 11716
rect 18095 11713 18107 11714
rect 18049 11707 18107 11713
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 15948 11648 16865 11676
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 17052 11676 17080 11707
rect 17218 11676 17224 11688
rect 17052 11648 17224 11676
rect 16853 11639 16911 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 17368 11648 17461 11676
rect 17368 11636 17374 11648
rect 18136 11645 18153 11676
rect 18187 11645 18199 11679
rect 18414 11676 18420 11688
rect 18375 11648 18420 11676
rect 18136 11639 18199 11645
rect 14516 11580 14964 11608
rect 14516 11568 14522 11580
rect 16390 11568 16396 11620
rect 16448 11608 16454 11620
rect 17328 11608 17356 11636
rect 16448 11580 17356 11608
rect 18136 11608 18164 11639
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 19168 11676 19196 11716
rect 19306 11704 19340 11716
rect 19392 11744 19398 11756
rect 19720 11747 19748 11784
rect 19794 11747 19800 11756
rect 19392 11716 19656 11744
rect 19720 11719 19800 11747
rect 19392 11704 19398 11716
rect 19306 11676 19334 11704
rect 19168 11648 19334 11676
rect 19628 11676 19656 11716
rect 19794 11704 19800 11719
rect 19852 11744 19858 11756
rect 20070 11744 20076 11756
rect 19852 11716 19897 11744
rect 20031 11716 20076 11744
rect 19852 11704 19858 11716
rect 20070 11704 20076 11716
rect 20128 11704 20134 11756
rect 20898 11744 20904 11756
rect 20180 11716 20904 11744
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 19628 11648 19901 11676
rect 19889 11645 19901 11648
rect 19935 11645 19947 11679
rect 19889 11639 19947 11645
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11676 20039 11679
rect 20180 11676 20208 11716
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 21174 11744 21180 11756
rect 21135 11716 21180 11744
rect 21174 11704 21180 11716
rect 21232 11704 21238 11756
rect 21468 11753 21496 11852
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 22005 11883 22063 11889
rect 22005 11880 22017 11883
rect 21968 11852 22017 11880
rect 21968 11840 21974 11852
rect 22005 11849 22017 11852
rect 22051 11849 22063 11883
rect 22005 11843 22063 11849
rect 21542 11772 21548 11824
rect 21600 11812 21606 11824
rect 22157 11815 22215 11821
rect 22157 11812 22169 11815
rect 21600 11784 22169 11812
rect 21600 11772 21606 11784
rect 22157 11781 22169 11784
rect 22203 11781 22215 11815
rect 22157 11775 22215 11781
rect 22373 11815 22431 11821
rect 22373 11781 22385 11815
rect 22419 11812 22431 11815
rect 22738 11812 22744 11824
rect 22419 11784 22744 11812
rect 22419 11781 22431 11784
rect 22373 11775 22431 11781
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 22388 11744 22416 11775
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 21499 11716 22416 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 20027 11648 20208 11676
rect 20027 11645 20039 11648
rect 19981 11639 20039 11645
rect 19150 11608 19156 11620
rect 18136 11580 19156 11608
rect 16448 11568 16454 11580
rect 19150 11568 19156 11580
rect 19208 11608 19214 11620
rect 19996 11608 20024 11639
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 21284 11676 21312 11707
rect 37366 11704 37372 11756
rect 37424 11744 37430 11756
rect 37461 11747 37519 11753
rect 37461 11744 37473 11747
rect 37424 11716 37473 11744
rect 37424 11704 37430 11716
rect 37461 11713 37473 11716
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 20312 11648 22232 11676
rect 20312 11636 20318 11648
rect 21450 11608 21456 11620
rect 19208 11580 20024 11608
rect 21411 11580 21456 11608
rect 19208 11568 19214 11580
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 16206 11540 16212 11552
rect 13004 11512 16212 11540
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 16356 11512 17233 11540
rect 16356 11500 16362 11512
rect 17221 11509 17233 11512
rect 17267 11540 17279 11543
rect 20162 11540 20168 11552
rect 17267 11512 20168 11540
rect 17267 11509 17279 11512
rect 17221 11503 17279 11509
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 21174 11500 21180 11552
rect 21232 11540 21238 11552
rect 21542 11540 21548 11552
rect 21232 11512 21548 11540
rect 21232 11500 21238 11512
rect 21542 11500 21548 11512
rect 21600 11500 21606 11552
rect 22204 11549 22232 11648
rect 22189 11543 22247 11549
rect 22189 11509 22201 11543
rect 22235 11509 22247 11543
rect 22189 11503 22247 11509
rect 37553 11543 37611 11549
rect 37553 11509 37565 11543
rect 37599 11540 37611 11543
rect 38102 11540 38108 11552
rect 37599 11512 38108 11540
rect 37599 11509 37611 11512
rect 37553 11503 37611 11509
rect 38102 11500 38108 11512
rect 38160 11500 38166 11552
rect 38286 11540 38292 11552
rect 38247 11512 38292 11540
rect 38286 11500 38292 11512
rect 38344 11500 38350 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 12250 11336 12256 11348
rect 12211 11308 12256 11336
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12618 11336 12624 11348
rect 12400 11308 12624 11336
rect 12400 11296 12406 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 12952 11308 14381 11336
rect 12952 11296 12958 11308
rect 14369 11305 14381 11308
rect 14415 11336 14427 11339
rect 15838 11336 15844 11348
rect 14415 11308 15844 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 18414 11336 18420 11348
rect 16040 11308 18420 11336
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 16040 11268 16068 11308
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 21174 11336 21180 11348
rect 20395 11308 21180 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 10560 11240 16068 11268
rect 16209 11271 16267 11277
rect 10560 11228 10566 11240
rect 16209 11237 16221 11271
rect 16255 11268 16267 11271
rect 17218 11268 17224 11280
rect 16255 11240 17224 11268
rect 16255 11237 16267 11240
rect 16209 11231 16267 11237
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 21818 11268 21824 11280
rect 18564 11240 21824 11268
rect 18564 11228 18570 11240
rect 21818 11228 21824 11240
rect 21876 11228 21882 11280
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 3050 11200 3056 11212
rect 3007 11172 3056 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 16025 11203 16083 11209
rect 11839 11172 12434 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 3476 11104 3521 11132
rect 3476 11092 3482 11104
rect 3234 11064 3240 11076
rect 3195 11036 3240 11064
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 12406 11064 12434 11172
rect 16025 11169 16037 11203
rect 16071 11200 16083 11203
rect 16390 11200 16396 11212
rect 16071 11172 16396 11200
rect 16071 11169 16083 11172
rect 16025 11163 16083 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 19794 11160 19800 11212
rect 19852 11200 19858 11212
rect 37182 11200 37188 11212
rect 19852 11172 20484 11200
rect 37143 11172 37188 11200
rect 19852 11160 19858 11172
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 14458 11132 14464 11144
rect 14419 11104 14464 11132
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 16298 11132 16304 11144
rect 16259 11104 16304 11132
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 20162 11092 20168 11144
rect 20220 11132 20226 11144
rect 20456 11141 20484 11172
rect 37182 11160 37188 11172
rect 37240 11160 37246 11212
rect 38102 11200 38108 11212
rect 38063 11172 38108 11200
rect 38102 11160 38108 11172
rect 38160 11160 38166 11212
rect 38286 11200 38292 11212
rect 38247 11172 38292 11200
rect 38286 11160 38292 11172
rect 38344 11160 38350 11212
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 20220 11104 20269 11132
rect 20220 11092 20226 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11101 20499 11135
rect 20441 11095 20499 11101
rect 18322 11064 18328 11076
rect 12406 11036 18328 11064
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 16264 10968 16313 10996
rect 16264 10956 16270 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 18340 10996 18368 11024
rect 20806 10996 20812 11008
rect 18340 10968 20812 10996
rect 16301 10959 16359 10965
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3234 10792 3240 10804
rect 2823 10764 3240 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 2958 10656 2964 10668
rect 2915 10628 2964 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18380 10628 18429 10656
rect 18380 10616 18386 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 3418 10588 3424 10600
rect 2179 10560 3424 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 18598 10588 18604 10600
rect 18559 10560 18604 10588
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 19426 10588 19432 10600
rect 19387 10560 19432 10588
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 18509 10251 18567 10257
rect 18509 10217 18521 10251
rect 18555 10248 18567 10251
rect 18598 10248 18604 10260
rect 18555 10220 18604 10248
rect 18555 10217 18567 10220
rect 18509 10211 18567 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 18414 10044 18420 10056
rect 18375 10016 18420 10044
rect 18414 10004 18420 10016
rect 18472 10044 18478 10056
rect 32950 10044 32956 10056
rect 18472 10016 32956 10044
rect 18472 10004 18478 10016
rect 32950 10004 32956 10016
rect 33008 10004 33014 10056
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2516 9500 2544 9531
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 23201 9571 23259 9577
rect 23201 9568 23213 9571
rect 2924 9540 23213 9568
rect 2924 9528 2930 9540
rect 23201 9537 23213 9540
rect 23247 9537 23259 9571
rect 23842 9568 23848 9580
rect 23803 9540 23848 9568
rect 23201 9531 23259 9537
rect 4706 9500 4712 9512
rect 2516 9472 4712 9500
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 23216 9432 23244 9531
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 23293 9503 23351 9509
rect 23293 9469 23305 9503
rect 23339 9500 23351 9503
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 23339 9472 24041 9500
rect 23339 9469 23351 9472
rect 23293 9463 23351 9469
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 25685 9503 25743 9509
rect 25685 9469 25697 9503
rect 25731 9500 25743 9503
rect 34514 9500 34520 9512
rect 25731 9472 34520 9500
rect 25731 9469 25743 9472
rect 25685 9463 25743 9469
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 29086 9432 29092 9444
rect 23216 9404 29092 9432
rect 29086 9392 29092 9404
rect 29144 9392 29150 9444
rect 2038 9364 2044 9376
rect 1999 9336 2044 9364
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 3234 9364 3240 9376
rect 2639 9336 3240 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2038 9052 2044 9104
rect 2096 9092 2102 9104
rect 2096 9064 3464 9092
rect 2096 9052 2102 9064
rect 3234 9024 3240 9036
rect 3195 8996 3240 9024
rect 3234 8984 3240 8996
rect 3292 8984 3298 9036
rect 3436 9033 3464 9064
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 8993 3479 9027
rect 3421 8987 3479 8993
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 34790 8956 34796 8968
rect 4764 8928 34796 8956
rect 4764 8916 4770 8928
rect 34790 8916 34796 8928
rect 34848 8916 34854 8968
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8956 37887 8959
rect 38286 8956 38292 8968
rect 37875 8928 38292 8956
rect 37875 8925 37887 8928
rect 37829 8919 37887 8925
rect 38286 8916 38292 8928
rect 38344 8916 38350 8968
rect 1578 8888 1584 8900
rect 1539 8860 1584 8888
rect 1578 8848 1584 8860
rect 1636 8848 1642 8900
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 20346 8480 20352 8492
rect 1903 8452 20352 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 37826 8276 37832 8288
rect 37787 8248 37832 8276
rect 37826 8236 37832 8248
rect 37884 8236 37890 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 37182 7936 37188 7948
rect 37143 7908 37188 7936
rect 37182 7896 37188 7908
rect 37240 7896 37246 7948
rect 37826 7896 37832 7948
rect 37884 7936 37890 7948
rect 38289 7939 38347 7945
rect 38289 7936 38301 7939
rect 37884 7908 38301 7936
rect 37884 7896 37890 7908
rect 38289 7905 38301 7908
rect 38335 7905 38347 7939
rect 38289 7899 38347 7905
rect 37550 7760 37556 7812
rect 37608 7800 37614 7812
rect 38105 7803 38163 7809
rect 38105 7800 38117 7803
rect 37608 7772 38117 7800
rect 37608 7760 37614 7772
rect 38105 7769 38117 7772
rect 38151 7769 38163 7803
rect 38105 7763 38163 7769
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 37550 7528 37556 7540
rect 37511 7500 37556 7528
rect 37550 7488 37556 7500
rect 37608 7488 37614 7540
rect 37366 7352 37372 7404
rect 37424 7392 37430 7404
rect 37461 7395 37519 7401
rect 37461 7392 37473 7395
rect 37424 7364 37473 7392
rect 37424 7352 37430 7364
rect 37461 7361 37473 7364
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 38010 7352 38016 7404
rect 38068 7392 38074 7404
rect 38105 7395 38163 7401
rect 38105 7392 38117 7395
rect 38068 7364 38117 7392
rect 38068 7352 38074 7364
rect 38105 7361 38117 7364
rect 38151 7361 38163 7395
rect 38105 7355 38163 7361
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 3418 7188 3424 7200
rect 2179 7160 3424 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 5350 7188 5356 7200
rect 5311 7160 5356 7188
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 38102 7148 38108 7200
rect 38160 7188 38166 7200
rect 38197 7191 38255 7197
rect 38197 7188 38209 7191
rect 38160 7160 38209 7188
rect 38160 7148 38166 7160
rect 38197 7157 38209 7160
rect 38243 7157 38255 7191
rect 38197 7151 38255 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3418 6848 3424 6860
rect 3379 6820 3424 6848
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 5350 6848 5356 6860
rect 5311 6820 5356 6848
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5810 6848 5816 6860
rect 5771 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 37182 6848 37188 6860
rect 37143 6820 37188 6848
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 38102 6848 38108 6860
rect 38063 6820 38108 6848
rect 38102 6808 38108 6820
rect 38160 6808 38166 6860
rect 38286 6848 38292 6860
rect 38247 6820 38292 6848
rect 38286 6808 38292 6820
rect 38344 6808 38350 6860
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 2464 6684 3249 6712
rect 2464 6672 2470 6684
rect 3237 6681 3249 6684
rect 3283 6681 3295 6715
rect 5534 6712 5540 6724
rect 5495 6684 5540 6712
rect 3237 6675 3295 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2406 6440 2412 6452
rect 2367 6412 2412 6440
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 4706 6372 4712 6384
rect 2516 6344 4712 6372
rect 2516 6316 2544 6344
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 4120 6276 5457 6304
rect 4120 6264 4126 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 37274 6264 37280 6316
rect 37332 6304 37338 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37332 6276 37473 6304
rect 37332 6264 37338 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 37553 6103 37611 6109
rect 37553 6069 37565 6103
rect 37599 6100 37611 6103
rect 38102 6100 38108 6112
rect 37599 6072 38108 6100
rect 37599 6069 37611 6072
rect 37553 6063 37611 6069
rect 38102 6060 38108 6072
rect 38160 6060 38166 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 39298 5828 39304 5840
rect 37844 5800 39304 5828
rect 37844 5769 37872 5800
rect 39298 5788 39304 5800
rect 39356 5788 39362 5840
rect 37829 5763 37887 5769
rect 37829 5729 37841 5763
rect 37875 5729 37887 5763
rect 38102 5760 38108 5772
rect 38063 5732 38108 5760
rect 37829 5723 37887 5729
rect 38102 5720 38108 5732
rect 38160 5720 38166 5772
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1912 5664 1961 5692
rect 1912 5652 1918 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 3142 5692 3148 5704
rect 2823 5664 3148 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3602 5692 3608 5704
rect 3283 5664 3608 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3602 5652 3608 5664
rect 3660 5692 3666 5704
rect 20806 5692 20812 5704
rect 3660 5664 20812 5692
rect 3660 5652 3666 5664
rect 20806 5652 20812 5664
rect 20864 5652 20870 5704
rect 38286 5652 38292 5704
rect 38344 5692 38350 5704
rect 38344 5664 38389 5692
rect 38344 5652 38350 5664
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3510 5556 3516 5568
rect 3375 5528 3516 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 37829 5219 37887 5225
rect 37829 5185 37841 5219
rect 37875 5216 37887 5219
rect 38286 5216 38292 5228
rect 37875 5188 38292 5216
rect 37875 5185 37887 5188
rect 37829 5179 37887 5185
rect 38286 5176 38292 5188
rect 38344 5176 38350 5228
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2222 5148 2228 5160
rect 2087 5120 2228 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2222 5108 2228 5120
rect 2280 5108 2286 5160
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 14 5040 20 5092
rect 72 5080 78 5092
rect 2332 5080 2360 5111
rect 72 5052 2360 5080
rect 72 5040 78 5052
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 4706 5012 4712 5024
rect 4203 4984 4712 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 36906 5012 36912 5024
rect 36867 4984 36912 5012
rect 36906 4972 36912 4984
rect 36964 4972 36970 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 2682 4672 2688 4684
rect 2332 4644 2688 4672
rect 2332 4613 2360 4644
rect 2682 4632 2688 4644
rect 2740 4672 2746 4684
rect 37090 4672 37096 4684
rect 2740 4644 5028 4672
rect 37051 4644 37096 4672
rect 2740 4632 2746 4644
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 2777 4567 2835 4573
rect 2792 4536 2820 4567
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 5000 4613 5028 4644
rect 37090 4632 37096 4644
rect 37148 4632 37154 4684
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 8294 4604 8300 4616
rect 8255 4576 8300 4604
rect 4985 4567 5043 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 25866 4564 25872 4616
rect 25924 4604 25930 4616
rect 25961 4607 26019 4613
rect 25961 4604 25973 4607
rect 25924 4576 25973 4604
rect 25924 4564 25930 4576
rect 25961 4573 25973 4576
rect 26007 4573 26019 4607
rect 25961 4567 26019 4573
rect 38194 4564 38200 4616
rect 38252 4604 38258 4616
rect 38252 4576 38297 4604
rect 38252 4564 38258 4576
rect 3326 4536 3332 4548
rect 2792 4508 3332 4536
rect 3326 4496 3332 4508
rect 3384 4536 3390 4548
rect 19334 4536 19340 4548
rect 3384 4508 19340 4536
rect 3384 4496 3390 4508
rect 19334 4496 19340 4508
rect 19392 4496 19398 4548
rect 38010 4536 38016 4548
rect 37971 4508 38016 4536
rect 38010 4496 38016 4508
rect 38068 4496 38074 4548
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3786 4468 3792 4480
rect 2915 4440 3792 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 5077 4471 5135 4477
rect 5077 4437 5089 4471
rect 5123 4468 5135 4471
rect 5718 4468 5724 4480
rect 5123 4440 5724 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3786 4196 3792 4208
rect 3747 4168 3792 4196
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 10502 4128 10508 4140
rect 10463 4100 10508 4128
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 24946 4128 24952 4140
rect 24907 4100 24952 4128
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 25961 4131 26019 4137
rect 25961 4097 25973 4131
rect 26007 4097 26019 4131
rect 37458 4128 37464 4140
rect 37419 4100 37464 4128
rect 25961 4091 26019 4097
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3200 4032 3985 4060
rect 3200 4020 3206 4032
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 3973 4023 4031 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8536 4032 8677 4060
rect 8536 4020 8542 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 25976 3992 26004 4091
rect 37458 4088 37464 4100
rect 37516 4088 37522 4140
rect 35802 4060 35808 4072
rect 35763 4032 35808 4060
rect 35802 4020 35808 4032
rect 35860 4020 35866 4072
rect 36725 4063 36783 4069
rect 36725 4029 36737 4063
rect 36771 4029 36783 4063
rect 36725 4023 36783 4029
rect 36909 4063 36967 4069
rect 36909 4029 36921 4063
rect 36955 4060 36967 4063
rect 38105 4063 38163 4069
rect 38105 4060 38117 4063
rect 36955 4032 38117 4060
rect 36955 4029 36967 4032
rect 36909 4023 36967 4029
rect 38105 4029 38117 4032
rect 38151 4029 38163 4063
rect 38105 4023 38163 4029
rect 2372 3964 26004 3992
rect 36740 3992 36768 4023
rect 37553 3995 37611 4001
rect 37553 3992 37565 3995
rect 36740 3964 37565 3992
rect 2372 3952 2378 3964
rect 37553 3961 37565 3964
rect 37599 3961 37611 3995
rect 37553 3955 37611 3961
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 4614 3924 4620 3936
rect 4479 3896 4620 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19484 3896 19625 3924
rect 19484 3884 19490 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 20714 3924 20720 3936
rect 20675 3896 20720 3924
rect 19613 3887 19671 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 22002 3924 22008 3936
rect 21963 3896 22008 3924
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 24854 3924 24860 3936
rect 24815 3896 24860 3924
rect 24854 3884 24860 3896
rect 24912 3884 24918 3936
rect 26050 3924 26056 3936
rect 26011 3896 26056 3924
rect 26050 3884 26056 3896
rect 26108 3884 26114 3936
rect 30006 3924 30012 3936
rect 29967 3896 30012 3924
rect 30006 3884 30012 3896
rect 30064 3884 30070 3936
rect 33962 3924 33968 3936
rect 33923 3896 33968 3924
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 34790 3884 34796 3936
rect 34848 3924 34854 3936
rect 37458 3924 37464 3936
rect 34848 3896 37464 3924
rect 34848 3884 34854 3896
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 5442 3720 5448 3732
rect 3936 3692 5448 3720
rect 3936 3680 3942 3692
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5626 3652 5632 3664
rect 5368 3624 5632 3652
rect 2774 3584 2780 3596
rect 2735 3556 2780 3584
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 3970 3584 3976 3596
rect 3467 3556 3976 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5368 3516 5396 3624
rect 5626 3612 5632 3624
rect 5684 3652 5690 3664
rect 10870 3652 10876 3664
rect 5684 3624 10876 3652
rect 5684 3612 5690 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 37366 3652 37372 3664
rect 28368 3624 37372 3652
rect 5534 3584 5540 3596
rect 5495 3556 5540 3584
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 10594 3584 10600 3596
rect 10555 3556 10600 3584
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 20714 3584 20720 3596
rect 20675 3556 20720 3584
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 25866 3584 25872 3596
rect 25827 3556 25872 3584
rect 25866 3544 25872 3556
rect 25924 3544 25930 3596
rect 26050 3584 26056 3596
rect 26011 3556 26056 3584
rect 26050 3544 26056 3556
rect 26108 3544 26114 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 5031 3488 5396 3516
rect 8573 3519 8631 3525
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8846 3516 8852 3528
rect 8619 3488 8852 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9766 3516 9772 3528
rect 9355 3488 9772 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9999 3488 10425 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12952 3488 13001 3516
rect 12952 3476 12958 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19392 3488 19625 3516
rect 19392 3476 19398 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3516 19763 3519
rect 19978 3516 19984 3528
rect 19751 3488 19984 3516
rect 19751 3485 19763 3488
rect 19705 3479 19763 3485
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 24302 3516 24308 3528
rect 23247 3488 24308 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 24302 3476 24308 3488
rect 24360 3476 24366 3528
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24636 3488 24685 3516
rect 24636 3476 24642 3488
rect 24673 3485 24685 3488
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 28258 3476 28264 3528
rect 28316 3516 28322 3528
rect 28368 3525 28396 3624
rect 37366 3612 37372 3624
rect 37424 3612 37430 3664
rect 29086 3544 29092 3596
rect 29144 3544 29150 3596
rect 30006 3584 30012 3596
rect 29967 3556 30012 3584
rect 30006 3544 30012 3556
rect 30064 3544 30070 3596
rect 35897 3587 35955 3593
rect 35897 3553 35909 3587
rect 35943 3584 35955 3587
rect 36262 3584 36268 3596
rect 35943 3556 36268 3584
rect 35943 3553 35955 3556
rect 35897 3547 35955 3553
rect 36262 3544 36268 3556
rect 36320 3544 36326 3596
rect 28353 3519 28411 3525
rect 28353 3516 28365 3519
rect 28316 3488 28365 3516
rect 28316 3476 28322 3488
rect 28353 3485 28365 3488
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 28997 3519 29055 3525
rect 28997 3485 29009 3519
rect 29043 3516 29055 3519
rect 29104 3516 29132 3544
rect 33870 3516 33876 3528
rect 29043 3488 29132 3516
rect 33831 3488 33876 3516
rect 29043 3485 29055 3488
rect 28997 3479 29055 3485
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35253 3519 35311 3525
rect 35253 3516 35265 3519
rect 34848 3488 35265 3516
rect 34848 3476 34854 3488
rect 35253 3485 35265 3488
rect 35299 3485 35311 3519
rect 35253 3479 35311 3485
rect 3234 3448 3240 3460
rect 3195 3420 3240 3448
rect 3234 3408 3240 3420
rect 3292 3408 3298 3460
rect 7377 3451 7435 3457
rect 7377 3417 7389 3451
rect 7423 3448 7435 3451
rect 20898 3448 20904 3460
rect 7423 3420 11928 3448
rect 7423 3417 7435 3420
rect 7377 3411 7435 3417
rect 4338 3340 4344 3392
rect 4396 3380 4402 3392
rect 4893 3383 4951 3389
rect 4893 3380 4905 3383
rect 4396 3352 4905 3380
rect 4396 3340 4402 3352
rect 4893 3349 4905 3352
rect 4939 3349 4951 3383
rect 4893 3343 4951 3349
rect 9030 3340 9036 3392
rect 9088 3380 9094 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 9088 3352 9229 3380
rect 9088 3340 9094 3352
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 11900 3380 11928 3420
rect 12406 3420 19840 3448
rect 20859 3420 20904 3448
rect 12406 3380 12434 3420
rect 11900 3352 12434 3380
rect 9217 3343 9275 3349
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 19518 3380 19524 3392
rect 19392 3352 19524 3380
rect 19392 3340 19398 3352
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 19812 3380 19840 3420
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 29089 3451 29147 3457
rect 29089 3417 29101 3451
rect 29135 3448 29147 3451
rect 30193 3451 30251 3457
rect 30193 3448 30205 3451
rect 29135 3420 30205 3448
rect 29135 3417 29147 3420
rect 29089 3411 29147 3417
rect 30193 3417 30205 3420
rect 30239 3417 30251 3451
rect 30193 3411 30251 3417
rect 31849 3451 31907 3457
rect 31849 3417 31861 3451
rect 31895 3448 31907 3451
rect 34054 3448 34060 3460
rect 31895 3420 34060 3448
rect 31895 3417 31907 3420
rect 31849 3411 31907 3417
rect 34054 3408 34060 3420
rect 34112 3408 34118 3460
rect 35345 3451 35403 3457
rect 35345 3417 35357 3451
rect 35391 3448 35403 3451
rect 36081 3451 36139 3457
rect 36081 3448 36093 3451
rect 35391 3420 36093 3448
rect 35391 3417 35403 3420
rect 35345 3411 35403 3417
rect 36081 3417 36093 3420
rect 36127 3417 36139 3451
rect 36081 3411 36139 3417
rect 37737 3451 37795 3457
rect 37737 3417 37749 3451
rect 37783 3448 37795 3451
rect 38654 3448 38660 3460
rect 37783 3420 38660 3448
rect 37783 3417 37795 3420
rect 37737 3411 37795 3417
rect 38654 3408 38660 3420
rect 38712 3408 38718 3460
rect 24394 3380 24400 3392
rect 19812 3352 24400 3380
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 28074 3340 28080 3392
rect 28132 3380 28138 3392
rect 28261 3383 28319 3389
rect 28261 3380 28273 3383
rect 28132 3352 28273 3380
rect 28132 3340 28138 3352
rect 28261 3349 28273 3352
rect 28307 3349 28319 3383
rect 28261 3343 28319 3349
rect 33965 3383 34023 3389
rect 33965 3349 33977 3383
rect 34011 3380 34023 3383
rect 34146 3380 34152 3392
rect 34011 3352 34152 3380
rect 34011 3349 34023 3352
rect 33965 3343 34023 3349
rect 34146 3340 34152 3352
rect 34204 3340 34210 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 658 3136 664 3188
rect 716 3176 722 3188
rect 37553 3179 37611 3185
rect 716 3148 5580 3176
rect 716 3136 722 3148
rect 3510 3108 3516 3120
rect 3471 3080 3516 3108
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 2866 2972 2872 2984
rect 2827 2944 2872 2972
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 4706 2972 4712 2984
rect 3743 2944 4712 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 3326 2864 3332 2916
rect 3384 2904 3390 2916
rect 4816 2904 4844 2935
rect 3384 2876 4844 2904
rect 5552 2904 5580 3148
rect 37553 3145 37565 3179
rect 37599 3176 37611 3179
rect 38010 3176 38016 3188
rect 37599 3148 38016 3176
rect 37599 3145 37611 3148
rect 37553 3139 37611 3145
rect 38010 3136 38016 3148
rect 38068 3136 38074 3188
rect 9030 3108 9036 3120
rect 8991 3080 9036 3108
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 19705 3111 19763 3117
rect 19705 3077 19717 3111
rect 19751 3108 19763 3111
rect 19978 3108 19984 3120
rect 19751 3080 19984 3108
rect 19751 3077 19763 3080
rect 19705 3071 19763 3077
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 28074 3108 28080 3120
rect 28035 3080 28080 3108
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 34146 3108 34152 3120
rect 34107 3080 34152 3108
rect 34146 3068 34152 3080
rect 34204 3068 34210 3120
rect 8846 3040 8852 3052
rect 8807 3012 8852 3040
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 11940 3012 12265 3040
rect 11940 3000 11946 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 12894 3040 12900 3052
rect 12855 3012 12900 3040
rect 12253 3003 12311 3009
rect 6546 2972 6552 2984
rect 6507 2944 6552 2972
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2972 6791 2975
rect 7466 2972 7472 2984
rect 6779 2944 7472 2972
rect 6779 2941 6791 2944
rect 6733 2935 6791 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 9309 2935 9367 2941
rect 9324 2904 9352 2935
rect 5552 2876 9352 2904
rect 12268 2904 12296 3003
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 19484 3012 19533 3040
rect 19484 3000 19490 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 19521 3003 19579 3009
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 24302 3040 24308 3052
rect 24263 3012 24308 3040
rect 24302 3000 24308 3012
rect 24360 3000 24366 3052
rect 33962 3040 33968 3052
rect 33923 3012 33968 3040
rect 33962 3000 33968 3012
rect 34020 3000 34026 3052
rect 36262 3040 36268 3052
rect 36223 3012 36268 3040
rect 36262 3000 36268 3012
rect 36320 3000 36326 3052
rect 37458 3040 37464 3052
rect 37419 3012 37464 3040
rect 37458 3000 37464 3012
rect 37516 3000 37522 3052
rect 38105 3043 38163 3049
rect 38105 3009 38117 3043
rect 38151 3040 38163 3043
rect 38194 3040 38200 3052
rect 38151 3012 38200 3040
rect 38151 3009 38163 3012
rect 38105 3003 38163 3009
rect 38194 3000 38200 3012
rect 38252 3000 38258 3052
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2972 12403 2975
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 12391 2944 13093 2972
rect 12391 2941 12403 2944
rect 12345 2935 12403 2941
rect 13081 2941 13093 2944
rect 13127 2941 13139 2975
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 13081 2935 13139 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 22186 2972 22192 2984
rect 22147 2944 22192 2972
rect 22186 2932 22192 2944
rect 22244 2932 22250 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24486 2972 24492 2984
rect 24447 2944 24492 2972
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 24765 2975 24823 2981
rect 24765 2941 24777 2975
rect 24811 2941 24823 2975
rect 27890 2972 27896 2984
rect 27851 2944 27896 2972
rect 24765 2935 24823 2941
rect 22002 2904 22008 2916
rect 12268 2876 22008 2904
rect 3384 2864 3390 2876
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 23198 2864 23204 2916
rect 23256 2904 23262 2916
rect 24780 2904 24808 2935
rect 27890 2932 27896 2944
rect 27948 2932 27954 2984
rect 28350 2972 28356 2984
rect 28311 2944 28356 2972
rect 28350 2932 28356 2944
rect 28408 2932 28414 2984
rect 34790 2972 34796 2984
rect 34751 2944 34796 2972
rect 34790 2932 34796 2944
rect 34848 2932 34854 2984
rect 23256 2876 24808 2904
rect 23256 2864 23262 2876
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 4706 2836 4712 2848
rect 2648 2808 4712 2836
rect 2648 2796 2654 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 3234 2632 3240 2644
rect 2547 2604 3240 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6604 2604 6745 2632
rect 6604 2592 6610 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 6733 2595 6791 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 8444 2604 8493 2632
rect 8444 2592 8450 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 14734 2632 14740 2644
rect 9815 2604 14740 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 20809 2635 20867 2641
rect 20809 2601 20821 2635
rect 20855 2632 20867 2635
rect 20898 2632 20904 2644
rect 20855 2604 20904 2632
rect 20855 2601 20867 2604
rect 20809 2595 20867 2601
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 22097 2635 22155 2641
rect 22097 2601 22109 2635
rect 22143 2632 22155 2635
rect 22186 2632 22192 2644
rect 22143 2604 22192 2632
rect 22143 2601 22155 2604
rect 22097 2595 22155 2601
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 23017 2635 23075 2641
rect 23017 2601 23029 2635
rect 23063 2632 23075 2635
rect 24486 2632 24492 2644
rect 23063 2604 24492 2632
rect 23063 2601 23075 2604
rect 23017 2595 23075 2601
rect 24486 2592 24492 2604
rect 24544 2592 24550 2644
rect 27890 2592 27896 2644
rect 27948 2632 27954 2644
rect 27985 2635 28043 2641
rect 27985 2632 27997 2635
rect 27948 2604 27997 2632
rect 27948 2592 27954 2604
rect 27985 2601 27997 2604
rect 28031 2601 28043 2635
rect 27985 2595 28043 2601
rect 4798 2564 4804 2576
rect 3252 2536 4804 2564
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2498 2388 2504 2440
rect 2556 2428 2562 2440
rect 3252 2437 3280 2536
rect 4798 2524 4804 2536
rect 4856 2564 4862 2576
rect 10321 2567 10379 2573
rect 4856 2536 6914 2564
rect 4856 2524 4862 2536
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 4614 2496 4620 2508
rect 4019 2468 4620 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 4764 2468 4809 2496
rect 4764 2456 4770 2468
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2556 2400 2605 2428
rect 2556 2388 2562 2400
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 6886 2428 6914 2536
rect 10321 2533 10333 2567
rect 10367 2533 10379 2567
rect 10321 2527 10379 2533
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 6886 2400 7573 2428
rect 3237 2391 3295 2397
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10336 2428 10364 2527
rect 10870 2524 10876 2576
rect 10928 2564 10934 2576
rect 10928 2536 12388 2564
rect 10928 2524 10934 2536
rect 10980 2437 11008 2536
rect 11790 2496 11796 2508
rect 11751 2468 11796 2496
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12250 2496 12256 2508
rect 12211 2468 12256 2496
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 12360 2496 12388 2536
rect 13998 2524 14004 2576
rect 14056 2564 14062 2576
rect 31021 2567 31079 2573
rect 31021 2564 31033 2567
rect 14056 2536 31033 2564
rect 14056 2524 14062 2536
rect 31021 2533 31033 2536
rect 31067 2533 31079 2567
rect 37182 2564 37188 2576
rect 31021 2527 31079 2533
rect 36464 2536 37188 2564
rect 17494 2496 17500 2508
rect 12360 2468 17500 2496
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 24578 2496 24584 2508
rect 24539 2468 24584 2496
rect 24578 2456 24584 2468
rect 24636 2456 24642 2508
rect 24765 2499 24823 2505
rect 24765 2465 24777 2499
rect 24811 2496 24823 2499
rect 24854 2496 24860 2508
rect 24811 2468 24860 2496
rect 24811 2465 24823 2468
rect 24765 2459 24823 2465
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 25130 2496 25136 2508
rect 25091 2468 25136 2496
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 29914 2456 29920 2508
rect 29972 2496 29978 2508
rect 36464 2505 36492 2536
rect 37182 2524 37188 2536
rect 37240 2524 37246 2576
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 29972 2468 30021 2496
rect 29972 2456 29978 2468
rect 30009 2465 30021 2468
rect 30055 2465 30067 2499
rect 30009 2459 30067 2465
rect 36449 2499 36507 2505
rect 36449 2465 36461 2499
rect 36495 2465 36507 2499
rect 36906 2496 36912 2508
rect 36867 2468 36912 2496
rect 36449 2459 36507 2465
rect 36906 2456 36912 2468
rect 36964 2456 36970 2508
rect 37642 2456 37648 2508
rect 37700 2456 37706 2508
rect 9907 2400 10364 2428
rect 10505 2431 10563 2437
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 20806 2428 20812 2440
rect 20763 2400 20812 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 3329 2363 3387 2369
rect 3329 2329 3341 2363
rect 3375 2360 3387 2363
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3375 2332 4169 2360
rect 3375 2329 3387 2332
rect 3329 2323 3387 2329
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 8588 2292 8616 2391
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 10520 2360 10548 2391
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 22002 2428 22008 2440
rect 21915 2400 22008 2428
rect 22002 2388 22008 2400
rect 22060 2428 22066 2440
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22060 2400 22937 2428
rect 22060 2388 22066 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29052 2400 29745 2428
rect 29052 2388 29058 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2428 37611 2431
rect 37660 2428 37688 2456
rect 37599 2400 37688 2428
rect 37599 2397 37611 2400
rect 37553 2391 37611 2397
rect 9088 2332 10548 2360
rect 11057 2363 11115 2369
rect 9088 2320 9094 2332
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11103 2332 11989 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 28258 2360 28264 2372
rect 17460 2332 28264 2360
rect 17460 2320 17466 2332
rect 28258 2320 28264 2332
rect 28316 2320 28322 2372
rect 30926 2320 30932 2372
rect 30984 2360 30990 2372
rect 31205 2363 31263 2369
rect 31205 2360 31217 2363
rect 30984 2332 31217 2360
rect 30984 2320 30990 2332
rect 31205 2329 31217 2332
rect 31251 2329 31263 2363
rect 31205 2323 31263 2329
rect 36725 2363 36783 2369
rect 36725 2329 36737 2363
rect 36771 2360 36783 2363
rect 37645 2363 37703 2369
rect 37645 2360 37657 2363
rect 36771 2332 37657 2360
rect 36771 2329 36783 2332
rect 36725 2323 36783 2329
rect 37645 2329 37657 2332
rect 37691 2329 37703 2363
rect 37645 2323 37703 2329
rect 9674 2292 9680 2304
rect 8588 2264 9680 2292
rect 9674 2252 9680 2264
rect 9732 2292 9738 2304
rect 17218 2292 17224 2304
rect 9732 2264 17224 2292
rect 9732 2252 9738 2264
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 17494 2252 17500 2304
rect 17552 2292 17558 2304
rect 24946 2292 24952 2304
rect 17552 2264 24952 2292
rect 17552 2252 17558 2264
rect 24946 2252 24952 2264
rect 25004 2252 25010 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 37832 37612 37884 37664
rect 39304 37612 39356 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2412 37272 2464 37324
rect 19156 37272 19208 37324
rect 25780 37315 25832 37324
rect 25780 37281 25789 37315
rect 25789 37281 25823 37315
rect 25823 37281 25832 37315
rect 25780 37272 25832 37281
rect 28632 37315 28684 37324
rect 28632 37281 28641 37315
rect 28641 37281 28675 37315
rect 28675 37281 28684 37315
rect 28632 37272 28684 37281
rect 30288 37272 30340 37324
rect 32864 37272 32916 37324
rect 33048 37272 33100 37324
rect 35348 37272 35400 37324
rect 38292 37315 38344 37324
rect 38292 37281 38301 37315
rect 38301 37281 38335 37315
rect 38335 37281 38344 37315
rect 38292 37272 38344 37281
rect 20 37204 72 37256
rect 2504 37247 2556 37256
rect 2504 37213 2513 37247
rect 2513 37213 2547 37247
rect 2547 37213 2556 37247
rect 2504 37204 2556 37213
rect 3424 37247 3476 37256
rect 3424 37213 3433 37247
rect 3433 37213 3467 37247
rect 3467 37213 3476 37247
rect 3424 37204 3476 37213
rect 4160 37247 4212 37256
rect 4160 37213 4169 37247
rect 4169 37213 4203 37247
rect 4203 37213 4212 37247
rect 4160 37204 4212 37213
rect 6552 37247 6604 37256
rect 6552 37213 6561 37247
rect 6561 37213 6595 37247
rect 6595 37213 6604 37247
rect 6552 37204 6604 37213
rect 9220 37247 9272 37256
rect 9220 37213 9229 37247
rect 9229 37213 9263 37247
rect 9263 37213 9272 37247
rect 9220 37204 9272 37213
rect 14464 37247 14516 37256
rect 14464 37213 14473 37247
rect 14473 37213 14507 37247
rect 14507 37213 14516 37247
rect 14464 37204 14516 37213
rect 14924 37247 14976 37256
rect 14924 37213 14933 37247
rect 14933 37213 14967 37247
rect 14967 37213 14976 37247
rect 14924 37204 14976 37213
rect 16212 37204 16264 37256
rect 17592 37247 17644 37256
rect 17592 37213 17601 37247
rect 17601 37213 17635 37247
rect 17635 37213 17644 37247
rect 17592 37204 17644 37213
rect 18880 37247 18932 37256
rect 18880 37213 18889 37247
rect 18889 37213 18923 37247
rect 18923 37213 18932 37247
rect 18880 37204 18932 37213
rect 19432 37204 19484 37256
rect 20996 37247 21048 37256
rect 20996 37213 21005 37247
rect 21005 37213 21039 37247
rect 21039 37213 21048 37247
rect 20996 37204 21048 37213
rect 22744 37247 22796 37256
rect 5356 37136 5408 37188
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 27804 37247 27856 37256
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 32496 37247 32548 37256
rect 26240 37136 26292 37188
rect 26424 37179 26476 37188
rect 26424 37145 26433 37179
rect 26433 37145 26467 37179
rect 26467 37145 26476 37179
rect 26424 37136 26476 37145
rect 4344 37068 4396 37120
rect 14648 37068 14700 37120
rect 18696 37068 18748 37120
rect 22284 37068 22336 37120
rect 32496 37213 32505 37247
rect 32505 37213 32539 37247
rect 32539 37213 32548 37247
rect 32496 37204 32548 37213
rect 36912 37247 36964 37256
rect 36912 37213 36921 37247
rect 36921 37213 36955 37247
rect 36955 37213 36964 37247
rect 38016 37247 38068 37256
rect 36912 37204 36964 37213
rect 38016 37213 38025 37247
rect 38025 37213 38059 37247
rect 38059 37213 38068 37247
rect 38016 37204 38068 37213
rect 30104 37179 30156 37188
rect 30104 37145 30113 37179
rect 30113 37145 30147 37179
rect 30147 37145 30156 37179
rect 30104 37136 30156 37145
rect 32680 37179 32732 37188
rect 32680 37145 32689 37179
rect 32689 37145 32723 37179
rect 32723 37145 32732 37179
rect 32680 37136 32732 37145
rect 30656 37068 30708 37120
rect 38200 37136 38252 37188
rect 38660 37068 38712 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 17592 36864 17644 36916
rect 23480 36864 23532 36916
rect 26240 36864 26292 36916
rect 38200 36907 38252 36916
rect 1860 36839 1912 36848
rect 1860 36805 1869 36839
rect 1869 36805 1903 36839
rect 1903 36805 1912 36839
rect 1860 36796 1912 36805
rect 2504 36796 2556 36848
rect 4344 36839 4396 36848
rect 4344 36805 4353 36839
rect 4353 36805 4387 36839
rect 4387 36805 4396 36839
rect 4344 36796 4396 36805
rect 14648 36839 14700 36848
rect 14648 36805 14657 36839
rect 14657 36805 14691 36839
rect 14691 36805 14700 36839
rect 14648 36796 14700 36805
rect 16764 36796 16816 36848
rect 22284 36839 22336 36848
rect 22284 36805 22293 36839
rect 22293 36805 22327 36839
rect 22327 36805 22336 36839
rect 22284 36796 22336 36805
rect 4160 36771 4212 36780
rect 4160 36737 4169 36771
rect 4169 36737 4203 36771
rect 4203 36737 4212 36771
rect 4160 36728 4212 36737
rect 6552 36771 6604 36780
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 9220 36771 9272 36780
rect 9220 36737 9229 36771
rect 9229 36737 9263 36771
rect 9263 36737 9272 36771
rect 9220 36728 9272 36737
rect 19156 36771 19208 36780
rect 19156 36737 19165 36771
rect 19165 36737 19199 36771
rect 19199 36737 19208 36771
rect 19156 36728 19208 36737
rect 19432 36728 19484 36780
rect 23572 36728 23624 36780
rect 27804 36796 27856 36848
rect 31760 36796 31812 36848
rect 38200 36873 38209 36907
rect 38209 36873 38243 36907
rect 38243 36873 38252 36907
rect 38200 36864 38252 36873
rect 37464 36796 37516 36848
rect 3516 36703 3568 36712
rect 3516 36669 3525 36703
rect 3525 36669 3559 36703
rect 3559 36669 3568 36703
rect 3516 36660 3568 36669
rect 3240 36592 3292 36644
rect 6460 36660 6512 36712
rect 7104 36703 7156 36712
rect 7104 36669 7113 36703
rect 7113 36669 7147 36703
rect 7147 36669 7156 36703
rect 7104 36660 7156 36669
rect 9404 36703 9456 36712
rect 9404 36669 9413 36703
rect 9413 36669 9447 36703
rect 9447 36669 9456 36703
rect 9404 36660 9456 36669
rect 9680 36703 9732 36712
rect 9680 36669 9689 36703
rect 9689 36669 9723 36703
rect 9723 36669 9732 36703
rect 9680 36660 9732 36669
rect 14924 36660 14976 36712
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 18972 36703 19024 36712
rect 18972 36669 18981 36703
rect 18981 36669 19015 36703
rect 19015 36669 19024 36703
rect 18972 36660 19024 36669
rect 19892 36660 19944 36712
rect 20628 36660 20680 36712
rect 22744 36660 22796 36712
rect 22836 36703 22888 36712
rect 22836 36669 22845 36703
rect 22845 36669 22879 36703
rect 22879 36669 22888 36703
rect 24584 36703 24636 36712
rect 22836 36660 22888 36669
rect 24584 36669 24593 36703
rect 24593 36669 24627 36703
rect 24627 36669 24636 36703
rect 24584 36660 24636 36669
rect 27344 36703 27396 36712
rect 23848 36592 23900 36644
rect 27344 36669 27353 36703
rect 27353 36669 27387 36703
rect 27387 36669 27396 36703
rect 27344 36660 27396 36669
rect 29644 36703 29696 36712
rect 26516 36592 26568 36644
rect 28448 36592 28500 36644
rect 29644 36669 29653 36703
rect 29653 36669 29687 36703
rect 29687 36669 29696 36703
rect 29644 36660 29696 36669
rect 29736 36660 29788 36712
rect 32312 36703 32364 36712
rect 32312 36669 32321 36703
rect 32321 36669 32355 36703
rect 32355 36669 32364 36703
rect 32312 36660 32364 36669
rect 34612 36703 34664 36712
rect 32220 36592 32272 36644
rect 34612 36669 34621 36703
rect 34621 36669 34655 36703
rect 34655 36669 34664 36703
rect 34612 36660 34664 36669
rect 34796 36703 34848 36712
rect 34796 36669 34805 36703
rect 34805 36669 34839 36703
rect 34839 36669 34848 36703
rect 34796 36660 34848 36669
rect 34888 36660 34940 36712
rect 37188 36524 37240 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 6460 36363 6512 36372
rect 6460 36329 6469 36363
rect 6469 36329 6503 36363
rect 6503 36329 6512 36363
rect 6460 36320 6512 36329
rect 9404 36363 9456 36372
rect 9404 36329 9413 36363
rect 9413 36329 9447 36363
rect 9447 36329 9456 36363
rect 9404 36320 9456 36329
rect 19892 36363 19944 36372
rect 19892 36329 19901 36363
rect 19901 36329 19935 36363
rect 19935 36329 19944 36363
rect 19892 36320 19944 36329
rect 24584 36320 24636 36372
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 3424 36184 3476 36236
rect 4160 36184 4212 36236
rect 14464 36184 14516 36236
rect 16120 36227 16172 36236
rect 16120 36193 16129 36227
rect 16129 36193 16163 36227
rect 16163 36193 16172 36227
rect 16120 36184 16172 36193
rect 17408 36227 17460 36236
rect 17408 36193 17417 36227
rect 17417 36193 17451 36227
rect 17451 36193 17460 36227
rect 17408 36184 17460 36193
rect 18696 36227 18748 36236
rect 18696 36193 18705 36227
rect 18705 36193 18739 36227
rect 18739 36193 18748 36227
rect 18696 36184 18748 36193
rect 18880 36227 18932 36236
rect 18880 36193 18889 36227
rect 18889 36193 18923 36227
rect 18923 36193 18932 36227
rect 18880 36184 18932 36193
rect 20996 36227 21048 36236
rect 20996 36193 21005 36227
rect 21005 36193 21039 36227
rect 21039 36193 21048 36227
rect 20996 36184 21048 36193
rect 22100 36227 22152 36236
rect 22100 36193 22109 36227
rect 22109 36193 22143 36227
rect 22143 36193 22152 36227
rect 22100 36184 22152 36193
rect 25136 36227 25188 36236
rect 25136 36193 25145 36227
rect 25145 36193 25179 36227
rect 25179 36193 25188 36227
rect 25136 36184 25188 36193
rect 27068 36184 27120 36236
rect 29000 36184 29052 36236
rect 30932 36184 30984 36236
rect 37372 36252 37424 36304
rect 37188 36227 37240 36236
rect 37188 36193 37197 36227
rect 37197 36193 37231 36227
rect 37231 36193 37240 36227
rect 37188 36184 37240 36193
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 6368 36159 6420 36168
rect 6368 36125 6377 36159
rect 6377 36125 6411 36159
rect 6411 36125 6420 36159
rect 6368 36116 6420 36125
rect 1768 36091 1820 36100
rect 1768 36057 1777 36091
rect 1777 36057 1811 36091
rect 1811 36057 1820 36091
rect 1768 36048 1820 36057
rect 4160 36091 4212 36100
rect 4160 36057 4169 36091
rect 4169 36057 4203 36091
rect 4203 36057 4212 36091
rect 4160 36048 4212 36057
rect 8484 35980 8536 36032
rect 19340 36116 19392 36168
rect 24584 36159 24636 36168
rect 14924 36091 14976 36100
rect 14924 36057 14933 36091
rect 14933 36057 14967 36091
rect 14967 36057 14976 36091
rect 14924 36048 14976 36057
rect 21180 36091 21232 36100
rect 21180 36057 21189 36091
rect 21189 36057 21223 36091
rect 21223 36057 21232 36091
rect 21180 36048 21232 36057
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 26884 36159 26936 36168
rect 26884 36125 26893 36159
rect 26893 36125 26927 36159
rect 26927 36125 26936 36159
rect 26884 36116 26936 36125
rect 29092 36116 29144 36168
rect 32036 36159 32088 36168
rect 32036 36125 32045 36159
rect 32045 36125 32079 36159
rect 32079 36125 32088 36159
rect 32036 36116 32088 36125
rect 37648 36159 37700 36168
rect 37648 36125 37657 36159
rect 37657 36125 37691 36159
rect 37691 36125 37700 36159
rect 37648 36116 37700 36125
rect 24768 36091 24820 36100
rect 24768 36057 24777 36091
rect 24777 36057 24811 36091
rect 24811 36057 24820 36091
rect 24768 36048 24820 36057
rect 26608 36048 26660 36100
rect 29920 36091 29972 36100
rect 29920 36057 29929 36091
rect 29929 36057 29963 36091
rect 29963 36057 29972 36091
rect 29920 36048 29972 36057
rect 32220 36091 32272 36100
rect 32220 36057 32229 36091
rect 32229 36057 32263 36091
rect 32263 36057 32272 36091
rect 32220 36048 32272 36057
rect 15200 35980 15252 36032
rect 23296 35980 23348 36032
rect 25044 35980 25096 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1768 35776 1820 35828
rect 3516 35776 3568 35828
rect 4160 35776 4212 35828
rect 14924 35776 14976 35828
rect 15200 35776 15252 35828
rect 18972 35776 19024 35828
rect 21180 35776 21232 35828
rect 24768 35776 24820 35828
rect 26424 35776 26476 35828
rect 29920 35776 29972 35828
rect 32220 35776 32272 35828
rect 23296 35708 23348 35760
rect 27344 35708 27396 35760
rect 27712 35708 27764 35760
rect 28632 35708 28684 35760
rect 1584 35640 1636 35692
rect 2596 35640 2648 35692
rect 3332 35640 3384 35692
rect 3792 35640 3844 35692
rect 6368 35640 6420 35692
rect 15200 35683 15252 35692
rect 15200 35649 15209 35683
rect 15209 35649 15243 35683
rect 15243 35649 15252 35683
rect 15200 35640 15252 35649
rect 16948 35640 17000 35692
rect 18880 35683 18932 35692
rect 18880 35649 18889 35683
rect 18889 35649 18923 35683
rect 18923 35649 18932 35683
rect 18880 35640 18932 35649
rect 20720 35640 20772 35692
rect 23480 35640 23532 35692
rect 24584 35640 24636 35692
rect 25044 35683 25096 35692
rect 25044 35649 25053 35683
rect 25053 35649 25087 35683
rect 25087 35649 25096 35683
rect 25044 35640 25096 35649
rect 25964 35683 26016 35692
rect 25964 35649 25973 35683
rect 25973 35649 26007 35683
rect 26007 35649 26016 35683
rect 25964 35640 26016 35649
rect 35348 35708 35400 35760
rect 30196 35640 30248 35692
rect 30564 35683 30616 35692
rect 30564 35649 30573 35683
rect 30573 35649 30607 35683
rect 30607 35649 30616 35683
rect 30564 35640 30616 35649
rect 32036 35640 32088 35692
rect 38200 35640 38252 35692
rect 15292 35572 15344 35624
rect 27988 35572 28040 35624
rect 33048 35615 33100 35624
rect 33048 35581 33057 35615
rect 33057 35581 33091 35615
rect 33091 35581 33100 35615
rect 33048 35572 33100 35581
rect 34704 35572 34756 35624
rect 35808 35572 35860 35624
rect 37924 35504 37976 35556
rect 17868 35436 17920 35488
rect 36728 35436 36780 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 16948 35275 17000 35284
rect 16948 35241 16957 35275
rect 16957 35241 16991 35275
rect 16991 35241 17000 35275
rect 16948 35232 17000 35241
rect 18696 35275 18748 35284
rect 18696 35241 18705 35275
rect 18705 35241 18739 35275
rect 18739 35241 18748 35275
rect 18696 35232 18748 35241
rect 18880 35232 18932 35284
rect 26608 35275 26660 35284
rect 15384 35164 15436 35216
rect 26608 35241 26617 35275
rect 26617 35241 26651 35275
rect 26651 35241 26660 35275
rect 26608 35232 26660 35241
rect 26884 35232 26936 35284
rect 27988 35275 28040 35284
rect 27988 35241 27997 35275
rect 27997 35241 28031 35275
rect 28031 35241 28040 35275
rect 27988 35232 28040 35241
rect 29644 35232 29696 35284
rect 30104 35275 30156 35284
rect 30104 35241 30113 35275
rect 30113 35241 30147 35275
rect 30147 35241 30156 35275
rect 30104 35232 30156 35241
rect 30656 35275 30708 35284
rect 30656 35241 30665 35275
rect 30665 35241 30699 35275
rect 30699 35241 30708 35275
rect 30656 35232 30708 35241
rect 31760 35275 31812 35284
rect 31760 35241 31769 35275
rect 31769 35241 31803 35275
rect 31803 35241 31812 35275
rect 31760 35232 31812 35241
rect 32312 35275 32364 35284
rect 32312 35241 32321 35275
rect 32321 35241 32355 35275
rect 32355 35241 32364 35275
rect 32312 35232 32364 35241
rect 32680 35232 32732 35284
rect 34612 35232 34664 35284
rect 34796 35232 34848 35284
rect 35808 35232 35860 35284
rect 15292 35028 15344 35080
rect 17592 35028 17644 35080
rect 19432 35028 19484 35080
rect 20996 35028 21048 35080
rect 21272 35071 21324 35080
rect 21272 35037 21281 35071
rect 21281 35037 21315 35071
rect 21315 35037 21324 35071
rect 21272 35028 21324 35037
rect 25044 35096 25096 35148
rect 23388 35028 23440 35080
rect 26516 35071 26568 35080
rect 26516 35037 26525 35071
rect 26525 35037 26559 35071
rect 26559 35037 26568 35071
rect 26516 35028 26568 35037
rect 14648 34960 14700 35012
rect 18788 34960 18840 35012
rect 18880 35003 18932 35012
rect 18880 34969 18889 35003
rect 18889 34969 18923 35003
rect 18923 34969 18932 35003
rect 18880 34960 18932 34969
rect 15660 34935 15712 34944
rect 15660 34901 15669 34935
rect 15669 34901 15703 34935
rect 15703 34901 15712 34935
rect 15660 34892 15712 34901
rect 18144 34892 18196 34944
rect 19984 34935 20036 34944
rect 19984 34901 19993 34935
rect 19993 34901 20027 34935
rect 20027 34901 20036 34935
rect 19984 34892 20036 34901
rect 30196 35164 30248 35216
rect 33692 35164 33744 35216
rect 32312 34960 32364 35012
rect 33600 35028 33652 35080
rect 38200 35164 38252 35216
rect 37648 35096 37700 35148
rect 37832 35139 37884 35148
rect 37832 35105 37841 35139
rect 37841 35105 37875 35139
rect 37875 35105 37884 35139
rect 37832 35096 37884 35105
rect 22376 34892 22428 34944
rect 25412 34892 25464 34944
rect 25964 34892 26016 34944
rect 38292 35071 38344 35080
rect 38292 35037 38301 35071
rect 38301 35037 38335 35071
rect 38335 35037 38344 35071
rect 38292 35028 38344 35037
rect 37280 34960 37332 35012
rect 37556 34960 37608 35012
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2596 34688 2648 34740
rect 14832 34688 14884 34740
rect 15936 34688 15988 34740
rect 17592 34731 17644 34740
rect 17592 34697 17601 34731
rect 17601 34697 17635 34731
rect 17635 34697 17644 34731
rect 17592 34688 17644 34697
rect 19340 34688 19392 34740
rect 20996 34731 21048 34740
rect 20996 34697 21005 34731
rect 21005 34697 21039 34731
rect 21039 34697 21048 34731
rect 20996 34688 21048 34697
rect 30564 34688 30616 34740
rect 37556 34731 37608 34740
rect 18420 34620 18472 34672
rect 18880 34620 18932 34672
rect 22376 34620 22428 34672
rect 36728 34663 36780 34672
rect 36728 34629 36737 34663
rect 36737 34629 36771 34663
rect 36771 34629 36780 34663
rect 36728 34620 36780 34629
rect 37556 34697 37565 34731
rect 37565 34697 37599 34731
rect 37599 34697 37608 34731
rect 37556 34688 37608 34697
rect 37924 34620 37976 34672
rect 2412 34552 2464 34604
rect 3148 34552 3200 34604
rect 3332 34527 3384 34536
rect 3332 34493 3341 34527
rect 3341 34493 3375 34527
rect 3375 34493 3384 34527
rect 15384 34552 15436 34604
rect 18144 34595 18196 34604
rect 18144 34561 18153 34595
rect 18153 34561 18187 34595
rect 18187 34561 18196 34595
rect 18144 34552 18196 34561
rect 3332 34484 3384 34493
rect 15108 34484 15160 34536
rect 17408 34484 17460 34536
rect 17868 34484 17920 34536
rect 19984 34552 20036 34604
rect 22928 34595 22980 34604
rect 22928 34561 22937 34595
rect 22937 34561 22971 34595
rect 22971 34561 22980 34595
rect 22928 34552 22980 34561
rect 33600 34552 33652 34604
rect 37464 34595 37516 34604
rect 37464 34561 37473 34595
rect 37473 34561 37507 34595
rect 37507 34561 37516 34595
rect 37464 34552 37516 34561
rect 38292 34595 38344 34604
rect 38292 34561 38301 34595
rect 38301 34561 38335 34595
rect 38335 34561 38344 34595
rect 38292 34552 38344 34561
rect 18972 34484 19024 34536
rect 14740 34416 14792 34468
rect 20076 34484 20128 34536
rect 23756 34527 23808 34536
rect 23756 34493 23765 34527
rect 23765 34493 23799 34527
rect 23799 34493 23808 34527
rect 23756 34484 23808 34493
rect 24492 34527 24544 34536
rect 24492 34493 24501 34527
rect 24501 34493 24535 34527
rect 24535 34493 24544 34527
rect 24492 34484 24544 34493
rect 35716 34527 35768 34536
rect 35716 34493 35725 34527
rect 35725 34493 35759 34527
rect 35759 34493 35768 34527
rect 35716 34484 35768 34493
rect 37648 34484 37700 34536
rect 28448 34459 28500 34468
rect 14464 34391 14516 34400
rect 14464 34357 14473 34391
rect 14473 34357 14507 34391
rect 14507 34357 14516 34391
rect 14464 34348 14516 34357
rect 18696 34348 18748 34400
rect 28448 34425 28457 34459
rect 28457 34425 28491 34459
rect 28491 34425 28500 34459
rect 28448 34416 28500 34425
rect 29092 34459 29144 34468
rect 29092 34425 29101 34459
rect 29101 34425 29135 34459
rect 29135 34425 29144 34459
rect 29092 34416 29144 34425
rect 32496 34416 32548 34468
rect 20168 34348 20220 34400
rect 33784 34391 33836 34400
rect 33784 34357 33793 34391
rect 33793 34357 33827 34391
rect 33827 34357 33836 34391
rect 33784 34348 33836 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14648 34187 14700 34196
rect 14648 34153 14657 34187
rect 14657 34153 14691 34187
rect 14691 34153 14700 34187
rect 14648 34144 14700 34153
rect 18144 34144 18196 34196
rect 18420 34187 18472 34196
rect 18420 34153 18429 34187
rect 18429 34153 18463 34187
rect 18463 34153 18472 34187
rect 18420 34144 18472 34153
rect 20168 34144 20220 34196
rect 23388 34187 23440 34196
rect 23388 34153 23397 34187
rect 23397 34153 23431 34187
rect 23431 34153 23440 34187
rect 23388 34144 23440 34153
rect 15660 34008 15712 34060
rect 34704 34144 34756 34196
rect 36912 34144 36964 34196
rect 26976 34051 27028 34060
rect 26976 34017 26985 34051
rect 26985 34017 27019 34051
rect 27019 34017 27028 34051
rect 26976 34008 27028 34017
rect 33876 34008 33928 34060
rect 35440 34008 35492 34060
rect 38292 34051 38344 34060
rect 38292 34017 38301 34051
rect 38301 34017 38335 34051
rect 38335 34017 38344 34051
rect 38292 34008 38344 34017
rect 1860 33940 1912 33992
rect 3792 33940 3844 33992
rect 14464 33983 14516 33992
rect 14464 33949 14473 33983
rect 14473 33949 14507 33983
rect 14507 33949 14516 33983
rect 14464 33940 14516 33949
rect 16856 33983 16908 33992
rect 15108 33872 15160 33924
rect 16856 33949 16865 33983
rect 16865 33949 16899 33983
rect 16899 33949 16908 33983
rect 16856 33940 16908 33949
rect 17960 33940 18012 33992
rect 18696 33940 18748 33992
rect 18788 33940 18840 33992
rect 19248 33940 19300 33992
rect 21456 33983 21508 33992
rect 21456 33949 21465 33983
rect 21465 33949 21499 33983
rect 21499 33949 21508 33983
rect 21456 33940 21508 33949
rect 20996 33872 21048 33924
rect 21272 33872 21324 33924
rect 22468 33940 22520 33992
rect 25964 33983 26016 33992
rect 25964 33949 25973 33983
rect 25973 33949 26007 33983
rect 26007 33949 26016 33983
rect 25964 33940 26016 33949
rect 26792 33940 26844 33992
rect 27252 33940 27304 33992
rect 27896 33940 27948 33992
rect 36452 33983 36504 33992
rect 25504 33872 25556 33924
rect 36452 33949 36461 33983
rect 36461 33949 36495 33983
rect 36495 33949 36504 33983
rect 36452 33940 36504 33949
rect 32404 33915 32456 33924
rect 32404 33881 32413 33915
rect 32413 33881 32447 33915
rect 32447 33881 32456 33915
rect 32404 33872 32456 33881
rect 36820 33872 36872 33924
rect 2044 33804 2096 33856
rect 16580 33804 16632 33856
rect 18512 33804 18564 33856
rect 18880 33804 18932 33856
rect 21088 33804 21140 33856
rect 22836 33847 22888 33856
rect 22836 33813 22845 33847
rect 22845 33813 22879 33847
rect 22879 33813 22888 33847
rect 22836 33804 22888 33813
rect 24676 33804 24728 33856
rect 27160 33804 27212 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 16856 33600 16908 33652
rect 19248 33600 19300 33652
rect 21272 33643 21324 33652
rect 21272 33609 21281 33643
rect 21281 33609 21315 33643
rect 21315 33609 21324 33643
rect 21272 33600 21324 33609
rect 23756 33643 23808 33652
rect 23756 33609 23765 33643
rect 23765 33609 23799 33643
rect 23799 33609 23808 33643
rect 23756 33600 23808 33609
rect 25504 33643 25556 33652
rect 25504 33609 25513 33643
rect 25513 33609 25547 33643
rect 25547 33609 25556 33643
rect 25504 33600 25556 33609
rect 27252 33643 27304 33652
rect 27252 33609 27261 33643
rect 27261 33609 27295 33643
rect 27295 33609 27304 33643
rect 27252 33600 27304 33609
rect 32404 33643 32456 33652
rect 32404 33609 32413 33643
rect 32413 33609 32447 33643
rect 32447 33609 32456 33643
rect 32404 33600 32456 33609
rect 35348 33600 35400 33652
rect 36820 33643 36872 33652
rect 36820 33609 36829 33643
rect 36829 33609 36863 33643
rect 36863 33609 36872 33643
rect 36820 33600 36872 33609
rect 2044 33575 2096 33584
rect 2044 33541 2053 33575
rect 2053 33541 2087 33575
rect 2087 33541 2096 33575
rect 2044 33532 2096 33541
rect 17960 33532 18012 33584
rect 18604 33532 18656 33584
rect 24492 33575 24544 33584
rect 24492 33541 24501 33575
rect 24501 33541 24535 33575
rect 24535 33541 24544 33575
rect 24492 33532 24544 33541
rect 25596 33532 25648 33584
rect 33784 33575 33836 33584
rect 33784 33541 33793 33575
rect 33793 33541 33827 33575
rect 33827 33541 33836 33575
rect 33784 33532 33836 33541
rect 36452 33532 36504 33584
rect 1860 33507 1912 33516
rect 1860 33473 1869 33507
rect 1869 33473 1903 33507
rect 1903 33473 1912 33507
rect 1860 33464 1912 33473
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 15108 33507 15160 33516
rect 15108 33473 15117 33507
rect 15117 33473 15151 33507
rect 15151 33473 15160 33507
rect 15108 33464 15160 33473
rect 18144 33464 18196 33516
rect 19892 33507 19944 33516
rect 19892 33473 19901 33507
rect 19901 33473 19935 33507
rect 19935 33473 19944 33507
rect 19892 33464 19944 33473
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 2780 33396 2832 33405
rect 14740 33396 14792 33448
rect 18052 33396 18104 33448
rect 18972 33396 19024 33448
rect 20076 33507 20128 33516
rect 20076 33473 20085 33507
rect 20085 33473 20119 33507
rect 20119 33473 20128 33507
rect 21088 33507 21140 33516
rect 20076 33464 20128 33473
rect 21088 33473 21097 33507
rect 21097 33473 21131 33507
rect 21131 33473 21140 33507
rect 21088 33464 21140 33473
rect 23664 33507 23716 33516
rect 23664 33473 23673 33507
rect 23673 33473 23707 33507
rect 23707 33473 23716 33507
rect 23664 33464 23716 33473
rect 21272 33396 21324 33448
rect 20260 33371 20312 33380
rect 20260 33337 20269 33371
rect 20269 33337 20303 33371
rect 20303 33337 20312 33371
rect 20260 33328 20312 33337
rect 23664 33328 23716 33380
rect 26976 33464 27028 33516
rect 26792 33396 26844 33448
rect 27988 33464 28040 33516
rect 32312 33507 32364 33516
rect 32312 33473 32321 33507
rect 32321 33473 32355 33507
rect 32355 33473 32364 33507
rect 32312 33464 32364 33473
rect 33876 33396 33928 33448
rect 34520 33439 34572 33448
rect 34520 33405 34529 33439
rect 34529 33405 34563 33439
rect 34563 33405 34572 33439
rect 34520 33396 34572 33405
rect 37464 33464 37516 33516
rect 37372 33396 37424 33448
rect 14832 33303 14884 33312
rect 14832 33269 14841 33303
rect 14841 33269 14875 33303
rect 14875 33269 14884 33303
rect 14832 33260 14884 33269
rect 19984 33260 20036 33312
rect 20628 33260 20680 33312
rect 21364 33260 21416 33312
rect 24584 33260 24636 33312
rect 36360 33328 36412 33380
rect 28172 33260 28224 33312
rect 36452 33260 36504 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 20996 33099 21048 33108
rect 3884 32852 3936 32904
rect 10416 32895 10468 32904
rect 10416 32861 10425 32895
rect 10425 32861 10459 32895
rect 10459 32861 10468 32895
rect 10416 32852 10468 32861
rect 10600 32895 10652 32904
rect 10600 32861 10609 32895
rect 10609 32861 10643 32895
rect 10643 32861 10652 32895
rect 10600 32852 10652 32861
rect 14188 32852 14240 32904
rect 15200 32852 15252 32904
rect 14648 32827 14700 32836
rect 14648 32793 14682 32827
rect 14682 32793 14700 32827
rect 14648 32784 14700 32793
rect 16580 32827 16632 32836
rect 16580 32793 16614 32827
rect 16614 32793 16632 32827
rect 16580 32784 16632 32793
rect 16764 32784 16816 32836
rect 10508 32759 10560 32768
rect 10508 32725 10517 32759
rect 10517 32725 10551 32759
rect 10551 32725 10560 32759
rect 10508 32716 10560 32725
rect 12716 32759 12768 32768
rect 12716 32725 12725 32759
rect 12725 32725 12759 32759
rect 12759 32725 12768 32759
rect 12716 32716 12768 32725
rect 14924 32716 14976 32768
rect 17592 32716 17644 32768
rect 18788 32852 18840 32904
rect 20076 32988 20128 33040
rect 19984 32852 20036 32904
rect 20352 32895 20404 32904
rect 20352 32861 20361 32895
rect 20361 32861 20395 32895
rect 20395 32861 20404 32895
rect 20352 32852 20404 32861
rect 20996 33065 21005 33099
rect 21005 33065 21039 33099
rect 21039 33065 21048 33099
rect 20996 33056 21048 33065
rect 27068 33056 27120 33108
rect 21364 32988 21416 33040
rect 21272 32963 21324 32972
rect 21272 32929 21281 32963
rect 21281 32929 21315 32963
rect 21315 32929 21324 32963
rect 21272 32920 21324 32929
rect 21180 32895 21232 32904
rect 21180 32861 21189 32895
rect 21189 32861 21223 32895
rect 21223 32861 21232 32895
rect 21180 32852 21232 32861
rect 21364 32895 21416 32904
rect 21364 32861 21373 32895
rect 21373 32861 21407 32895
rect 21407 32861 21416 32895
rect 22376 32895 22428 32904
rect 21364 32852 21416 32861
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 22836 32852 22888 32904
rect 24952 32963 25004 32972
rect 24952 32929 24961 32963
rect 24961 32929 24995 32963
rect 24995 32929 25004 32963
rect 24952 32920 25004 32929
rect 25596 32988 25648 33040
rect 26700 32988 26752 33040
rect 26884 32920 26936 32972
rect 26056 32895 26108 32904
rect 18604 32784 18656 32836
rect 18696 32784 18748 32836
rect 19984 32759 20036 32768
rect 19984 32725 19993 32759
rect 19993 32725 20027 32759
rect 20027 32725 20036 32759
rect 19984 32716 20036 32725
rect 22468 32784 22520 32836
rect 24768 32827 24820 32836
rect 24768 32793 24777 32827
rect 24777 32793 24811 32827
rect 24811 32793 24820 32827
rect 24768 32784 24820 32793
rect 25136 32827 25188 32836
rect 25136 32793 25145 32827
rect 25145 32793 25179 32827
rect 25179 32793 25188 32827
rect 25136 32784 25188 32793
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 26240 32852 26292 32904
rect 26976 32852 27028 32904
rect 27344 32852 27396 32904
rect 27436 32895 27488 32904
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27896 32895 27948 32904
rect 27436 32852 27488 32861
rect 27896 32861 27905 32895
rect 27905 32861 27939 32895
rect 27939 32861 27948 32895
rect 27896 32852 27948 32861
rect 28172 32963 28224 32972
rect 28172 32929 28181 32963
rect 28181 32929 28215 32963
rect 28215 32929 28224 32963
rect 28172 32920 28224 32929
rect 28264 32895 28316 32904
rect 28264 32861 28273 32895
rect 28273 32861 28307 32895
rect 28307 32861 28316 32895
rect 28264 32852 28316 32861
rect 36452 32963 36504 32972
rect 36452 32929 36461 32963
rect 36461 32929 36495 32963
rect 36495 32929 36504 32963
rect 36452 32920 36504 32929
rect 38292 32963 38344 32972
rect 38292 32929 38301 32963
rect 38301 32929 38335 32963
rect 38335 32929 38344 32963
rect 38292 32920 38344 32929
rect 29000 32784 29052 32836
rect 36636 32827 36688 32836
rect 36636 32793 36645 32827
rect 36645 32793 36679 32827
rect 36679 32793 36688 32827
rect 36636 32784 36688 32793
rect 26608 32716 26660 32768
rect 27160 32716 27212 32768
rect 27528 32716 27580 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 14648 32555 14700 32564
rect 14648 32521 14657 32555
rect 14657 32521 14691 32555
rect 14691 32521 14700 32555
rect 14648 32512 14700 32521
rect 24492 32512 24544 32564
rect 26056 32512 26108 32564
rect 36636 32512 36688 32564
rect 2504 32444 2556 32496
rect 3884 32419 3936 32428
rect 3884 32385 3893 32419
rect 3893 32385 3927 32419
rect 3927 32385 3936 32419
rect 3884 32376 3936 32385
rect 10508 32376 10560 32428
rect 12716 32376 12768 32428
rect 14832 32419 14884 32428
rect 14832 32385 14841 32419
rect 14841 32385 14875 32419
rect 14875 32385 14884 32419
rect 14832 32376 14884 32385
rect 15016 32376 15068 32428
rect 16028 32376 16080 32428
rect 17408 32419 17460 32428
rect 17408 32385 17417 32419
rect 17417 32385 17451 32419
rect 17451 32385 17460 32419
rect 17408 32376 17460 32385
rect 17592 32419 17644 32428
rect 17592 32385 17601 32419
rect 17601 32385 17635 32419
rect 17635 32385 17644 32419
rect 17592 32376 17644 32385
rect 18512 32419 18564 32428
rect 18512 32385 18521 32419
rect 18521 32385 18555 32419
rect 18555 32385 18564 32419
rect 18512 32376 18564 32385
rect 18604 32376 18656 32428
rect 19432 32419 19484 32428
rect 2688 32351 2740 32360
rect 2688 32317 2697 32351
rect 2697 32317 2731 32351
rect 2731 32317 2740 32351
rect 2688 32308 2740 32317
rect 3700 32351 3752 32360
rect 3700 32317 3709 32351
rect 3709 32317 3743 32351
rect 3743 32317 3752 32351
rect 3700 32308 3752 32317
rect 8944 32308 8996 32360
rect 9404 32240 9456 32292
rect 12164 32351 12216 32360
rect 12164 32317 12173 32351
rect 12173 32317 12207 32351
rect 12207 32317 12216 32351
rect 12164 32308 12216 32317
rect 19156 32308 19208 32360
rect 19432 32385 19441 32419
rect 19441 32385 19475 32419
rect 19475 32385 19484 32419
rect 19432 32376 19484 32385
rect 20812 32376 20864 32428
rect 24676 32376 24728 32428
rect 26608 32376 26660 32428
rect 19984 32308 20036 32360
rect 20260 32308 20312 32360
rect 21364 32308 21416 32360
rect 9680 32172 9732 32224
rect 9956 32172 10008 32224
rect 20536 32240 20588 32292
rect 22468 32308 22520 32360
rect 25228 32351 25280 32360
rect 13544 32215 13596 32224
rect 13544 32181 13553 32215
rect 13553 32181 13587 32215
rect 13587 32181 13596 32215
rect 13544 32172 13596 32181
rect 15108 32172 15160 32224
rect 17316 32172 17368 32224
rect 18788 32172 18840 32224
rect 19616 32215 19668 32224
rect 19616 32181 19625 32215
rect 19625 32181 19659 32215
rect 19659 32181 19668 32215
rect 19616 32172 19668 32181
rect 25228 32317 25237 32351
rect 25237 32317 25271 32351
rect 25271 32317 25280 32351
rect 25228 32308 25280 32317
rect 25320 32351 25372 32360
rect 25320 32317 25329 32351
rect 25329 32317 25363 32351
rect 25363 32317 25372 32351
rect 25320 32308 25372 32317
rect 25504 32240 25556 32292
rect 26884 32444 26936 32496
rect 28540 32444 28592 32496
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 27252 32419 27304 32428
rect 27252 32385 27261 32419
rect 27261 32385 27295 32419
rect 27295 32385 27304 32419
rect 27528 32419 27580 32428
rect 27252 32376 27304 32385
rect 27528 32385 27537 32419
rect 27537 32385 27571 32419
rect 27571 32385 27580 32419
rect 27528 32376 27580 32385
rect 30564 32444 30616 32496
rect 29000 32419 29052 32428
rect 27068 32308 27120 32360
rect 29000 32385 29009 32419
rect 29009 32385 29043 32419
rect 29043 32385 29052 32419
rect 29000 32376 29052 32385
rect 36452 32419 36504 32428
rect 36452 32385 36461 32419
rect 36461 32385 36495 32419
rect 36495 32385 36504 32419
rect 36452 32376 36504 32385
rect 37648 32419 37700 32428
rect 37648 32385 37657 32419
rect 37657 32385 37691 32419
rect 37691 32385 37700 32419
rect 37648 32376 37700 32385
rect 29092 32351 29144 32360
rect 29092 32317 29101 32351
rect 29101 32317 29135 32351
rect 29135 32317 29144 32351
rect 29092 32308 29144 32317
rect 25044 32172 25096 32224
rect 27988 32240 28040 32292
rect 28724 32240 28776 32292
rect 31116 32172 31168 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 10416 32011 10468 32020
rect 10416 31977 10425 32011
rect 10425 31977 10459 32011
rect 10459 31977 10468 32011
rect 10416 31968 10468 31977
rect 12164 31968 12216 32020
rect 19616 32011 19668 32020
rect 4804 31900 4856 31952
rect 8944 31832 8996 31884
rect 1584 31764 1636 31816
rect 2504 31807 2556 31816
rect 2504 31773 2513 31807
rect 2513 31773 2547 31807
rect 2547 31773 2556 31807
rect 2504 31764 2556 31773
rect 9956 31764 10008 31816
rect 11796 31832 11848 31884
rect 19616 31977 19625 32011
rect 19625 31977 19659 32011
rect 19659 31977 19668 32011
rect 19616 31968 19668 31977
rect 19800 31968 19852 32020
rect 20628 31968 20680 32020
rect 24860 31968 24912 32020
rect 25320 31968 25372 32020
rect 27068 32011 27120 32020
rect 27068 31977 27077 32011
rect 27077 31977 27111 32011
rect 27111 31977 27120 32011
rect 27068 31968 27120 31977
rect 27988 31968 28040 32020
rect 28540 32011 28592 32020
rect 28540 31977 28549 32011
rect 28549 31977 28583 32011
rect 28583 31977 28592 32011
rect 28540 31968 28592 31977
rect 31116 32011 31168 32020
rect 31116 31977 31125 32011
rect 31125 31977 31159 32011
rect 31159 31977 31168 32011
rect 31116 31968 31168 31977
rect 13912 31900 13964 31952
rect 14924 31900 14976 31952
rect 15200 31832 15252 31884
rect 16028 31832 16080 31884
rect 9404 31739 9456 31748
rect 9404 31705 9413 31739
rect 9413 31705 9447 31739
rect 9447 31705 9456 31739
rect 9404 31696 9456 31705
rect 1768 31628 1820 31680
rect 9312 31671 9364 31680
rect 9312 31637 9321 31671
rect 9321 31637 9355 31671
rect 9355 31637 9364 31671
rect 9312 31628 9364 31637
rect 14280 31764 14332 31816
rect 13544 31696 13596 31748
rect 16672 31764 16724 31816
rect 17592 31764 17644 31816
rect 18328 31764 18380 31816
rect 20260 31832 20312 31884
rect 20536 31875 20588 31884
rect 20536 31841 20545 31875
rect 20545 31841 20579 31875
rect 20579 31841 20588 31875
rect 20536 31832 20588 31841
rect 20628 31875 20680 31884
rect 20628 31841 20637 31875
rect 20637 31841 20671 31875
rect 20671 31841 20680 31875
rect 20628 31832 20680 31841
rect 20996 31832 21048 31884
rect 18144 31739 18196 31748
rect 18144 31705 18153 31739
rect 18153 31705 18187 31739
rect 18187 31705 18196 31739
rect 18144 31696 18196 31705
rect 15384 31628 15436 31680
rect 15660 31628 15712 31680
rect 18420 31628 18472 31680
rect 19800 31807 19852 31816
rect 19800 31773 19809 31807
rect 19809 31773 19843 31807
rect 19843 31773 19852 31807
rect 19800 31764 19852 31773
rect 20076 31696 20128 31748
rect 19340 31628 19392 31680
rect 20812 31764 20864 31816
rect 22468 31900 22520 31952
rect 21456 31875 21508 31884
rect 21456 31841 21465 31875
rect 21465 31841 21499 31875
rect 21499 31841 21508 31875
rect 21456 31832 21508 31841
rect 25228 31900 25280 31952
rect 26976 31875 27028 31884
rect 20536 31696 20588 31748
rect 26976 31841 26985 31875
rect 26985 31841 27019 31875
rect 27019 31841 27028 31875
rect 26976 31832 27028 31841
rect 27804 31832 27856 31884
rect 25504 31764 25556 31816
rect 28264 31764 28316 31816
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 29736 31807 29788 31816
rect 29736 31773 29745 31807
rect 29745 31773 29779 31807
rect 29779 31773 29788 31807
rect 29736 31764 29788 31773
rect 33784 31807 33836 31816
rect 33784 31773 33793 31807
rect 33793 31773 33827 31807
rect 33827 31773 33836 31807
rect 33784 31764 33836 31773
rect 24400 31628 24452 31680
rect 27528 31696 27580 31748
rect 28080 31739 28132 31748
rect 28080 31705 28089 31739
rect 28089 31705 28123 31739
rect 28123 31705 28132 31739
rect 28080 31696 28132 31705
rect 30104 31696 30156 31748
rect 24768 31671 24820 31680
rect 24768 31637 24793 31671
rect 24793 31637 24820 31671
rect 24768 31628 24820 31637
rect 34060 31628 34112 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 3700 31424 3752 31476
rect 14188 31424 14240 31476
rect 18144 31467 18196 31476
rect 18144 31433 18153 31467
rect 18153 31433 18187 31467
rect 18187 31433 18196 31467
rect 18144 31424 18196 31433
rect 24952 31424 25004 31476
rect 25136 31467 25188 31476
rect 25136 31433 25145 31467
rect 25145 31433 25179 31467
rect 25179 31433 25188 31467
rect 25136 31424 25188 31433
rect 26240 31467 26292 31476
rect 26240 31433 26249 31467
rect 26249 31433 26283 31467
rect 26283 31433 26292 31467
rect 26240 31424 26292 31433
rect 28080 31424 28132 31476
rect 30104 31467 30156 31476
rect 30104 31433 30113 31467
rect 30113 31433 30147 31467
rect 30147 31433 30156 31467
rect 30104 31424 30156 31433
rect 2320 31331 2372 31340
rect 2320 31297 2329 31331
rect 2329 31297 2363 31331
rect 2363 31297 2372 31331
rect 2320 31288 2372 31297
rect 3608 31331 3660 31340
rect 3608 31297 3617 31331
rect 3617 31297 3651 31331
rect 3651 31297 3660 31331
rect 3608 31288 3660 31297
rect 9036 31288 9088 31340
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9723 31331
rect 9723 31297 9732 31331
rect 9680 31288 9732 31297
rect 15108 31288 15160 31340
rect 15844 31331 15896 31340
rect 15844 31297 15853 31331
rect 15853 31297 15887 31331
rect 15887 31297 15896 31331
rect 16028 31331 16080 31340
rect 15844 31288 15896 31297
rect 16028 31297 16037 31331
rect 16037 31297 16071 31331
rect 16071 31297 16080 31331
rect 16028 31288 16080 31297
rect 20720 31356 20772 31408
rect 24860 31356 24912 31408
rect 26148 31356 26200 31408
rect 27252 31356 27304 31408
rect 34060 31399 34112 31408
rect 34060 31365 34069 31399
rect 34069 31365 34103 31399
rect 34103 31365 34112 31399
rect 34060 31356 34112 31365
rect 35716 31399 35768 31408
rect 35716 31365 35725 31399
rect 35725 31365 35759 31399
rect 35759 31365 35768 31399
rect 35716 31356 35768 31365
rect 18420 31331 18472 31340
rect 18420 31297 18429 31331
rect 18429 31297 18463 31331
rect 18463 31297 18472 31331
rect 18420 31288 18472 31297
rect 24400 31331 24452 31340
rect 24400 31297 24409 31331
rect 24409 31297 24443 31331
rect 24443 31297 24452 31331
rect 24400 31288 24452 31297
rect 8576 31263 8628 31272
rect 8576 31229 8585 31263
rect 8585 31229 8619 31263
rect 8619 31229 8628 31263
rect 8576 31220 8628 31229
rect 9312 31220 9364 31272
rect 11060 31220 11112 31272
rect 11704 31220 11756 31272
rect 17224 31220 17276 31272
rect 18052 31220 18104 31272
rect 18328 31263 18380 31272
rect 18328 31229 18337 31263
rect 18337 31229 18371 31263
rect 18371 31229 18380 31263
rect 18328 31220 18380 31229
rect 21180 31220 21232 31272
rect 24676 31288 24728 31340
rect 25044 31331 25096 31340
rect 25044 31297 25053 31331
rect 25053 31297 25087 31331
rect 25087 31297 25096 31331
rect 25044 31288 25096 31297
rect 25596 31288 25648 31340
rect 25872 31331 25924 31340
rect 25872 31297 25881 31331
rect 25881 31297 25915 31331
rect 25915 31297 25924 31331
rect 25872 31288 25924 31297
rect 26240 31288 26292 31340
rect 26976 31288 27028 31340
rect 28172 31220 28224 31272
rect 28908 31220 28960 31272
rect 30564 31288 30616 31340
rect 33876 31263 33928 31272
rect 33876 31229 33885 31263
rect 33885 31229 33919 31263
rect 33919 31229 33928 31263
rect 33876 31220 33928 31229
rect 3240 31152 3292 31204
rect 8944 31195 8996 31204
rect 8944 31161 8953 31195
rect 8953 31161 8987 31195
rect 8987 31161 8996 31195
rect 8944 31152 8996 31161
rect 15292 31152 15344 31204
rect 26700 31152 26752 31204
rect 27344 31152 27396 31204
rect 2964 31127 3016 31136
rect 2964 31093 2973 31127
rect 2973 31093 3007 31127
rect 3007 31093 3016 31127
rect 2964 31084 3016 31093
rect 4068 31127 4120 31136
rect 4068 31093 4077 31127
rect 4077 31093 4111 31127
rect 4111 31093 4120 31127
rect 4068 31084 4120 31093
rect 9036 31127 9088 31136
rect 9036 31093 9045 31127
rect 9045 31093 9079 31127
rect 9079 31093 9088 31127
rect 9036 31084 9088 31093
rect 9496 31127 9548 31136
rect 9496 31093 9505 31127
rect 9505 31093 9539 31127
rect 9539 31093 9548 31127
rect 9496 31084 9548 31093
rect 14740 31084 14792 31136
rect 15016 31084 15068 31136
rect 19432 31084 19484 31136
rect 20536 31084 20588 31136
rect 38292 31084 38344 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3608 30880 3660 30932
rect 14280 30923 14332 30932
rect 14280 30889 14289 30923
rect 14289 30889 14323 30923
rect 14323 30889 14332 30923
rect 14280 30880 14332 30889
rect 15844 30880 15896 30932
rect 17224 30880 17276 30932
rect 15292 30812 15344 30864
rect 1584 30787 1636 30796
rect 1584 30753 1593 30787
rect 1593 30753 1627 30787
rect 1627 30753 1636 30787
rect 1584 30744 1636 30753
rect 1768 30787 1820 30796
rect 1768 30753 1777 30787
rect 1777 30753 1811 30787
rect 1811 30753 1820 30787
rect 1768 30744 1820 30753
rect 2780 30787 2832 30796
rect 2780 30753 2789 30787
rect 2789 30753 2823 30787
rect 2823 30753 2832 30787
rect 2780 30744 2832 30753
rect 9312 30744 9364 30796
rect 10140 30676 10192 30728
rect 11060 30719 11112 30728
rect 11060 30685 11069 30719
rect 11069 30685 11103 30719
rect 11103 30685 11112 30719
rect 11060 30676 11112 30685
rect 13360 30676 13412 30728
rect 14280 30744 14332 30796
rect 15016 30744 15068 30796
rect 15200 30744 15252 30796
rect 20628 30812 20680 30864
rect 25044 30880 25096 30932
rect 25596 30923 25648 30932
rect 25596 30889 25605 30923
rect 25605 30889 25639 30923
rect 25639 30889 25648 30923
rect 25596 30880 25648 30889
rect 26516 30880 26568 30932
rect 28264 30880 28316 30932
rect 28908 30880 28960 30932
rect 26700 30812 26752 30864
rect 18696 30744 18748 30796
rect 19064 30744 19116 30796
rect 17316 30676 17368 30728
rect 17960 30719 18012 30728
rect 17960 30685 17969 30719
rect 17969 30685 18003 30719
rect 18003 30685 18012 30719
rect 17960 30676 18012 30685
rect 18328 30676 18380 30728
rect 17408 30651 17460 30660
rect 2872 30540 2924 30592
rect 17408 30617 17417 30651
rect 17417 30617 17451 30651
rect 17451 30617 17460 30651
rect 17408 30608 17460 30617
rect 19340 30676 19392 30728
rect 20444 30744 20496 30796
rect 25872 30787 25924 30796
rect 25872 30753 25881 30787
rect 25881 30753 25915 30787
rect 25915 30753 25924 30787
rect 25872 30744 25924 30753
rect 26148 30744 26200 30796
rect 37832 30787 37884 30796
rect 37832 30753 37841 30787
rect 37841 30753 37875 30787
rect 37875 30753 37884 30787
rect 37832 30744 37884 30753
rect 38292 30787 38344 30796
rect 38292 30753 38301 30787
rect 38301 30753 38335 30787
rect 38335 30753 38344 30787
rect 38292 30744 38344 30753
rect 20076 30676 20128 30728
rect 22100 30719 22152 30728
rect 22100 30685 22109 30719
rect 22109 30685 22143 30719
rect 22143 30685 22152 30719
rect 22100 30676 22152 30685
rect 22376 30651 22428 30660
rect 22376 30617 22385 30651
rect 22385 30617 22419 30651
rect 22419 30617 22428 30651
rect 22376 30608 22428 30617
rect 26792 30676 26844 30728
rect 27252 30676 27304 30728
rect 27620 30719 27672 30728
rect 27620 30685 27629 30719
rect 27629 30685 27663 30719
rect 27663 30685 27672 30719
rect 27620 30676 27672 30685
rect 26240 30608 26292 30660
rect 28632 30608 28684 30660
rect 38108 30651 38160 30660
rect 38108 30617 38117 30651
rect 38117 30617 38151 30651
rect 38151 30617 38160 30651
rect 38108 30608 38160 30617
rect 13728 30583 13780 30592
rect 13728 30549 13737 30583
rect 13737 30549 13771 30583
rect 13771 30549 13780 30583
rect 13728 30540 13780 30549
rect 18236 30540 18288 30592
rect 18696 30583 18748 30592
rect 18696 30549 18705 30583
rect 18705 30549 18739 30583
rect 18739 30549 18748 30583
rect 18696 30540 18748 30549
rect 23112 30540 23164 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 15200 30379 15252 30388
rect 15200 30345 15209 30379
rect 15209 30345 15243 30379
rect 15243 30345 15252 30379
rect 15200 30336 15252 30345
rect 15844 30336 15896 30388
rect 17316 30379 17368 30388
rect 17316 30345 17325 30379
rect 17325 30345 17359 30379
rect 17359 30345 17368 30379
rect 17316 30336 17368 30345
rect 17408 30336 17460 30388
rect 23388 30336 23440 30388
rect 26516 30336 26568 30388
rect 27712 30336 27764 30388
rect 29736 30336 29788 30388
rect 38108 30336 38160 30388
rect 3148 30200 3200 30252
rect 4068 30243 4120 30252
rect 4068 30209 4077 30243
rect 4077 30209 4111 30243
rect 4111 30209 4120 30243
rect 4068 30200 4120 30209
rect 8576 30200 8628 30252
rect 9588 30268 9640 30320
rect 13728 30268 13780 30320
rect 15660 30268 15712 30320
rect 16028 30268 16080 30320
rect 16672 30268 16724 30320
rect 10140 30243 10192 30252
rect 10140 30209 10149 30243
rect 10149 30209 10183 30243
rect 10183 30209 10192 30243
rect 10140 30200 10192 30209
rect 11980 30200 12032 30252
rect 4620 30132 4672 30184
rect 3056 30064 3108 30116
rect 9496 30132 9548 30184
rect 9956 30132 10008 30184
rect 12164 30243 12216 30252
rect 12164 30209 12173 30243
rect 12173 30209 12207 30243
rect 12207 30209 12216 30243
rect 12164 30200 12216 30209
rect 13084 30200 13136 30252
rect 13544 30200 13596 30252
rect 14464 30200 14516 30252
rect 17960 30268 18012 30320
rect 18328 30311 18380 30320
rect 18328 30277 18337 30311
rect 18337 30277 18371 30311
rect 18371 30277 18380 30311
rect 18328 30268 18380 30277
rect 19432 30311 19484 30320
rect 19432 30277 19441 30311
rect 19441 30277 19475 30311
rect 19475 30277 19484 30311
rect 19432 30268 19484 30277
rect 19800 30268 19852 30320
rect 23112 30311 23164 30320
rect 19340 30200 19392 30252
rect 9404 30064 9456 30116
rect 2136 30039 2188 30048
rect 2136 30005 2145 30039
rect 2145 30005 2179 30039
rect 2179 30005 2188 30039
rect 2136 29996 2188 30005
rect 2872 30039 2924 30048
rect 2872 30005 2881 30039
rect 2881 30005 2915 30039
rect 2915 30005 2924 30039
rect 2872 29996 2924 30005
rect 7656 30039 7708 30048
rect 7656 30005 7665 30039
rect 7665 30005 7699 30039
rect 7699 30005 7708 30039
rect 7656 29996 7708 30005
rect 8944 29996 8996 30048
rect 11888 29996 11940 30048
rect 12164 30064 12216 30116
rect 17224 30132 17276 30184
rect 19156 30132 19208 30184
rect 20076 30200 20128 30252
rect 23112 30277 23121 30311
rect 23121 30277 23155 30311
rect 23155 30277 23164 30311
rect 23112 30268 23164 30277
rect 26056 30268 26108 30320
rect 30656 30311 30708 30320
rect 23020 30243 23072 30252
rect 23020 30209 23029 30243
rect 23029 30209 23063 30243
rect 23063 30209 23072 30243
rect 23020 30200 23072 30209
rect 23480 30200 23532 30252
rect 13912 30064 13964 30116
rect 15844 30064 15896 30116
rect 17500 30107 17552 30116
rect 13636 30039 13688 30048
rect 13636 30005 13645 30039
rect 13645 30005 13679 30039
rect 13679 30005 13688 30039
rect 13636 29996 13688 30005
rect 14924 29996 14976 30048
rect 15108 29996 15160 30048
rect 16948 30039 17000 30048
rect 16948 30005 16957 30039
rect 16957 30005 16991 30039
rect 16991 30005 17000 30039
rect 16948 29996 17000 30005
rect 17500 30073 17509 30107
rect 17509 30073 17543 30107
rect 17543 30073 17552 30107
rect 17500 30064 17552 30073
rect 17592 30064 17644 30116
rect 19892 30064 19944 30116
rect 19708 29996 19760 30048
rect 19984 29996 20036 30048
rect 22744 30132 22796 30184
rect 22376 30064 22428 30116
rect 24032 30200 24084 30252
rect 27804 30200 27856 30252
rect 28632 30200 28684 30252
rect 29828 30200 29880 30252
rect 30656 30277 30673 30311
rect 30673 30277 30708 30311
rect 30656 30268 30708 30277
rect 30012 30200 30064 30252
rect 31116 30200 31168 30252
rect 31576 30243 31628 30252
rect 31576 30209 31585 30243
rect 31585 30209 31619 30243
rect 31619 30209 31628 30243
rect 31576 30200 31628 30209
rect 32496 30200 32548 30252
rect 32680 30243 32732 30252
rect 32680 30209 32689 30243
rect 32689 30209 32723 30243
rect 32723 30209 32732 30243
rect 32680 30200 32732 30209
rect 37648 30200 37700 30252
rect 26516 30132 26568 30184
rect 24768 30064 24820 30116
rect 27528 30064 27580 30116
rect 27620 29996 27672 30048
rect 29000 29996 29052 30048
rect 29920 29996 29972 30048
rect 30932 30039 30984 30048
rect 30932 30005 30941 30039
rect 30941 30005 30975 30039
rect 30975 30005 30984 30039
rect 30932 29996 30984 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 4620 29792 4672 29844
rect 5356 29835 5408 29844
rect 5356 29801 5365 29835
rect 5365 29801 5399 29835
rect 5399 29801 5408 29835
rect 5356 29792 5408 29801
rect 10968 29792 11020 29844
rect 9128 29767 9180 29776
rect 9128 29733 9137 29767
rect 9137 29733 9171 29767
rect 9171 29733 9180 29767
rect 9128 29724 9180 29733
rect 11980 29792 12032 29844
rect 19800 29835 19852 29844
rect 14280 29767 14332 29776
rect 14280 29733 14289 29767
rect 14289 29733 14323 29767
rect 14323 29733 14332 29767
rect 14280 29724 14332 29733
rect 15292 29724 15344 29776
rect 17500 29724 17552 29776
rect 19800 29801 19809 29835
rect 19809 29801 19843 29835
rect 19843 29801 19852 29835
rect 19800 29792 19852 29801
rect 20628 29835 20680 29844
rect 20628 29801 20637 29835
rect 20637 29801 20671 29835
rect 20671 29801 20680 29835
rect 20628 29792 20680 29801
rect 22100 29792 22152 29844
rect 24860 29792 24912 29844
rect 26240 29792 26292 29844
rect 28632 29835 28684 29844
rect 28632 29801 28641 29835
rect 28641 29801 28675 29835
rect 28675 29801 28684 29835
rect 28632 29792 28684 29801
rect 29828 29792 29880 29844
rect 30564 29835 30616 29844
rect 30564 29801 30573 29835
rect 30573 29801 30607 29835
rect 30607 29801 30616 29835
rect 30564 29792 30616 29801
rect 33600 29792 33652 29844
rect 38384 29792 38436 29844
rect 2964 29656 3016 29708
rect 4620 29588 4672 29640
rect 1584 29563 1636 29572
rect 1584 29529 1593 29563
rect 1593 29529 1627 29563
rect 1627 29529 1636 29563
rect 1584 29520 1636 29529
rect 3240 29563 3292 29572
rect 3240 29529 3249 29563
rect 3249 29529 3283 29563
rect 3283 29529 3292 29563
rect 3240 29520 3292 29529
rect 10140 29656 10192 29708
rect 15660 29656 15712 29708
rect 7656 29588 7708 29640
rect 9588 29588 9640 29640
rect 10048 29631 10100 29640
rect 10048 29597 10057 29631
rect 10057 29597 10091 29631
rect 10091 29597 10100 29631
rect 10048 29588 10100 29597
rect 12440 29588 12492 29640
rect 2964 29452 3016 29504
rect 9036 29520 9088 29572
rect 11980 29520 12032 29572
rect 13636 29588 13688 29640
rect 14280 29588 14332 29640
rect 14464 29631 14516 29640
rect 14464 29597 14482 29631
rect 14482 29597 14516 29631
rect 14464 29588 14516 29597
rect 14740 29631 14792 29640
rect 14740 29597 14785 29631
rect 14785 29597 14792 29631
rect 14740 29588 14792 29597
rect 14924 29631 14976 29640
rect 14924 29597 14933 29631
rect 14933 29597 14967 29631
rect 14967 29597 14976 29631
rect 14924 29588 14976 29597
rect 15384 29588 15436 29640
rect 17132 29588 17184 29640
rect 17776 29588 17828 29640
rect 18604 29656 18656 29708
rect 23020 29656 23072 29708
rect 24676 29699 24728 29708
rect 24676 29665 24685 29699
rect 24685 29665 24719 29699
rect 24719 29665 24728 29699
rect 24676 29656 24728 29665
rect 26700 29699 26752 29708
rect 26700 29665 26709 29699
rect 26709 29665 26743 29699
rect 26743 29665 26752 29699
rect 26700 29656 26752 29665
rect 30932 29656 30984 29708
rect 37188 29699 37240 29708
rect 37188 29665 37197 29699
rect 37197 29665 37231 29699
rect 37231 29665 37240 29699
rect 37188 29656 37240 29665
rect 13360 29520 13412 29572
rect 12716 29452 12768 29504
rect 13268 29495 13320 29504
rect 13268 29461 13277 29495
rect 13277 29461 13311 29495
rect 13311 29461 13320 29495
rect 13268 29452 13320 29461
rect 13820 29452 13872 29504
rect 16856 29520 16908 29572
rect 18788 29520 18840 29572
rect 19524 29520 19576 29572
rect 19892 29588 19944 29640
rect 20076 29588 20128 29640
rect 20444 29588 20496 29640
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 20904 29588 20956 29640
rect 26516 29631 26568 29640
rect 26516 29597 26525 29631
rect 26525 29597 26559 29631
rect 26559 29597 26568 29631
rect 26516 29588 26568 29597
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 29920 29631 29972 29640
rect 29920 29597 29929 29631
rect 29929 29597 29963 29631
rect 29963 29597 29972 29631
rect 29920 29588 29972 29597
rect 31024 29588 31076 29640
rect 38292 29631 38344 29640
rect 38292 29597 38301 29631
rect 38301 29597 38335 29631
rect 38335 29597 38344 29631
rect 38292 29588 38344 29597
rect 23480 29520 23532 29572
rect 23756 29520 23808 29572
rect 27252 29563 27304 29572
rect 27252 29529 27261 29563
rect 27261 29529 27295 29563
rect 27295 29529 27304 29563
rect 27252 29520 27304 29529
rect 27896 29520 27948 29572
rect 29000 29520 29052 29572
rect 32312 29563 32364 29572
rect 32312 29529 32321 29563
rect 32321 29529 32355 29563
rect 32355 29529 32364 29563
rect 32312 29520 32364 29529
rect 32496 29563 32548 29572
rect 32496 29529 32505 29563
rect 32505 29529 32539 29563
rect 32539 29529 32548 29563
rect 32496 29520 32548 29529
rect 38108 29563 38160 29572
rect 38108 29529 38117 29563
rect 38117 29529 38151 29563
rect 38151 29529 38160 29563
rect 38108 29520 38160 29529
rect 15568 29452 15620 29504
rect 19432 29452 19484 29504
rect 20076 29452 20128 29504
rect 27344 29495 27396 29504
rect 27344 29461 27353 29495
rect 27353 29461 27387 29495
rect 27387 29461 27396 29495
rect 27344 29452 27396 29461
rect 29092 29452 29144 29504
rect 30656 29452 30708 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 10048 29248 10100 29300
rect 11888 29291 11940 29300
rect 11888 29257 11897 29291
rect 11897 29257 11931 29291
rect 11931 29257 11940 29291
rect 11888 29248 11940 29257
rect 12440 29248 12492 29300
rect 16764 29248 16816 29300
rect 16948 29248 17000 29300
rect 17224 29248 17276 29300
rect 2136 29155 2188 29164
rect 2136 29121 2145 29155
rect 2145 29121 2179 29155
rect 2179 29121 2188 29155
rect 2136 29112 2188 29121
rect 5356 29112 5408 29164
rect 2780 29044 2832 29096
rect 2872 29087 2924 29096
rect 2872 29053 2881 29087
rect 2881 29053 2915 29087
rect 2915 29053 2924 29087
rect 2872 29044 2924 29053
rect 4620 28976 4672 29028
rect 8668 29112 8720 29164
rect 10140 29112 10192 29164
rect 10968 29155 11020 29164
rect 10968 29121 10977 29155
rect 10977 29121 11011 29155
rect 11011 29121 11020 29155
rect 10968 29112 11020 29121
rect 11796 29112 11848 29164
rect 9680 29044 9732 29096
rect 12164 29044 12216 29096
rect 13820 29087 13872 29096
rect 13820 29053 13829 29087
rect 13829 29053 13863 29087
rect 13863 29053 13872 29087
rect 13820 29044 13872 29053
rect 14280 29044 14332 29096
rect 14740 29044 14792 29096
rect 15108 29112 15160 29164
rect 17132 29112 17184 29164
rect 18696 29180 18748 29232
rect 18788 29180 18840 29232
rect 24032 29180 24084 29232
rect 25964 29180 26016 29232
rect 32680 29248 32732 29300
rect 37648 29180 37700 29232
rect 15660 29044 15712 29096
rect 16948 29044 17000 29096
rect 21088 29112 21140 29164
rect 21180 29155 21232 29164
rect 21180 29121 21189 29155
rect 21189 29121 21223 29155
rect 21223 29121 21232 29155
rect 23388 29155 23440 29164
rect 21180 29112 21232 29121
rect 23388 29121 23397 29155
rect 23397 29121 23431 29155
rect 23431 29121 23440 29155
rect 23388 29112 23440 29121
rect 15292 28976 15344 29028
rect 15476 29019 15528 29028
rect 15476 28985 15485 29019
rect 15485 28985 15519 29019
rect 15519 28985 15528 29019
rect 15476 28976 15528 28985
rect 15568 29019 15620 29028
rect 15568 28985 15577 29019
rect 15577 28985 15611 29019
rect 15611 28985 15620 29019
rect 15568 28976 15620 28985
rect 15752 28976 15804 29028
rect 4712 28951 4764 28960
rect 4712 28917 4721 28951
rect 4721 28917 4755 28951
rect 4755 28917 4764 28951
rect 4712 28908 4764 28917
rect 7840 28951 7892 28960
rect 7840 28917 7849 28951
rect 7849 28917 7883 28951
rect 7883 28917 7892 28951
rect 7840 28908 7892 28917
rect 11888 28951 11940 28960
rect 11888 28917 11897 28951
rect 11897 28917 11931 28951
rect 11931 28917 11940 28951
rect 11888 28908 11940 28917
rect 13912 28908 13964 28960
rect 15384 28908 15436 28960
rect 25412 29044 25464 29096
rect 19156 28976 19208 29028
rect 26332 28976 26384 29028
rect 30012 29112 30064 29164
rect 31024 29112 31076 29164
rect 38292 29112 38344 29164
rect 30380 29087 30432 29096
rect 30380 29053 30389 29087
rect 30389 29053 30423 29087
rect 30423 29053 30432 29087
rect 30380 29044 30432 29053
rect 31576 29044 31628 29096
rect 18420 28908 18472 28960
rect 21180 28908 21232 28960
rect 26424 28908 26476 28960
rect 31392 28908 31444 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2780 28747 2832 28756
rect 2780 28713 2789 28747
rect 2789 28713 2823 28747
rect 2823 28713 2832 28747
rect 2780 28704 2832 28713
rect 11796 28747 11848 28756
rect 11796 28713 11805 28747
rect 11805 28713 11839 28747
rect 11839 28713 11848 28747
rect 11796 28704 11848 28713
rect 12164 28704 12216 28756
rect 16948 28747 17000 28756
rect 16948 28713 16957 28747
rect 16957 28713 16991 28747
rect 16991 28713 17000 28747
rect 16948 28704 17000 28713
rect 26516 28704 26568 28756
rect 28172 28747 28224 28756
rect 28172 28713 28181 28747
rect 28181 28713 28215 28747
rect 28215 28713 28224 28747
rect 28172 28704 28224 28713
rect 38108 28704 38160 28756
rect 20260 28636 20312 28688
rect 31576 28636 31628 28688
rect 4712 28568 4764 28620
rect 5632 28611 5684 28620
rect 5632 28577 5641 28611
rect 5641 28577 5675 28611
rect 5675 28577 5684 28611
rect 5632 28568 5684 28577
rect 7840 28568 7892 28620
rect 11888 28568 11940 28620
rect 17316 28568 17368 28620
rect 1860 28500 1912 28552
rect 2964 28500 3016 28552
rect 4252 28543 4304 28552
rect 4252 28509 4261 28543
rect 4261 28509 4295 28543
rect 4295 28509 4304 28543
rect 4252 28500 4304 28509
rect 9128 28500 9180 28552
rect 11980 28500 12032 28552
rect 17408 28500 17460 28552
rect 21272 28568 21324 28620
rect 27620 28568 27672 28620
rect 30012 28611 30064 28620
rect 30012 28577 30021 28611
rect 30021 28577 30055 28611
rect 30055 28577 30064 28611
rect 30012 28568 30064 28577
rect 37740 28568 37792 28620
rect 20812 28543 20864 28552
rect 20812 28509 20821 28543
rect 20821 28509 20855 28543
rect 20855 28509 20864 28543
rect 20812 28500 20864 28509
rect 20996 28500 21048 28552
rect 19156 28432 19208 28484
rect 20168 28432 20220 28484
rect 8760 28364 8812 28416
rect 11980 28407 12032 28416
rect 11980 28373 12007 28407
rect 12007 28373 12032 28407
rect 11980 28364 12032 28373
rect 20904 28364 20956 28416
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21824 28543 21876 28552
rect 21180 28500 21232 28509
rect 21824 28509 21833 28543
rect 21833 28509 21867 28543
rect 21867 28509 21876 28543
rect 21824 28500 21876 28509
rect 25228 28543 25280 28552
rect 25228 28509 25237 28543
rect 25237 28509 25271 28543
rect 25271 28509 25280 28543
rect 25228 28500 25280 28509
rect 28540 28500 28592 28552
rect 29000 28500 29052 28552
rect 30196 28500 30248 28552
rect 31392 28500 31444 28552
rect 35256 28500 35308 28552
rect 37924 28500 37976 28552
rect 23204 28407 23256 28416
rect 23204 28373 23213 28407
rect 23213 28373 23247 28407
rect 23247 28373 23256 28407
rect 23204 28364 23256 28373
rect 24400 28364 24452 28416
rect 25504 28475 25556 28484
rect 25504 28441 25538 28475
rect 25538 28441 25556 28475
rect 25504 28432 25556 28441
rect 30380 28432 30432 28484
rect 35992 28475 36044 28484
rect 35992 28441 36001 28475
rect 36001 28441 36035 28475
rect 36035 28441 36044 28475
rect 35992 28432 36044 28441
rect 37740 28432 37792 28484
rect 38200 28432 38252 28484
rect 26332 28364 26384 28416
rect 27804 28407 27856 28416
rect 27804 28373 27813 28407
rect 27813 28373 27847 28407
rect 27847 28373 27856 28407
rect 27804 28364 27856 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1860 28067 1912 28076
rect 1860 28033 1869 28067
rect 1869 28033 1903 28067
rect 1903 28033 1912 28067
rect 1860 28024 1912 28033
rect 4252 28024 4304 28076
rect 8852 28067 8904 28076
rect 8852 28033 8861 28067
rect 8861 28033 8895 28067
rect 8895 28033 8904 28067
rect 8852 28024 8904 28033
rect 11152 28024 11204 28076
rect 13268 28067 13320 28076
rect 13268 28033 13277 28067
rect 13277 28033 13311 28067
rect 13311 28033 13320 28067
rect 13268 28024 13320 28033
rect 2044 27999 2096 28008
rect 2044 27965 2053 27999
rect 2053 27965 2087 27999
rect 2087 27965 2096 27999
rect 2044 27956 2096 27965
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 2780 27956 2832 27965
rect 8760 27999 8812 28008
rect 8760 27965 8769 27999
rect 8769 27965 8803 27999
rect 8803 27965 8812 27999
rect 8760 27956 8812 27965
rect 11796 27999 11848 28008
rect 11796 27965 11805 27999
rect 11805 27965 11839 27999
rect 11839 27965 11848 27999
rect 11796 27956 11848 27965
rect 13360 27999 13412 28008
rect 13360 27965 13369 27999
rect 13369 27965 13403 27999
rect 13403 27965 13412 27999
rect 13360 27956 13412 27965
rect 15384 28024 15436 28076
rect 16212 28092 16264 28144
rect 19892 28160 19944 28212
rect 22928 28160 22980 28212
rect 24032 28160 24084 28212
rect 11060 27888 11112 27940
rect 15568 27956 15620 28008
rect 20260 28092 20312 28144
rect 23756 28135 23808 28144
rect 15752 27820 15804 27872
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 17684 27888 17736 27940
rect 20168 28024 20220 28076
rect 22744 28067 22796 28076
rect 22744 28033 22753 28067
rect 22753 28033 22787 28067
rect 22787 28033 22796 28067
rect 22744 28024 22796 28033
rect 23204 28024 23256 28076
rect 23756 28101 23765 28135
rect 23765 28101 23799 28135
rect 23799 28101 23808 28135
rect 23756 28092 23808 28101
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 26424 28160 26476 28212
rect 29092 28160 29144 28212
rect 32312 28203 32364 28212
rect 24400 28024 24452 28033
rect 20076 27956 20128 28008
rect 32312 28169 32321 28203
rect 32321 28169 32355 28203
rect 32355 28169 32364 28203
rect 32312 28160 32364 28169
rect 35256 28203 35308 28212
rect 35256 28169 35265 28203
rect 35265 28169 35299 28203
rect 35299 28169 35308 28203
rect 35256 28160 35308 28169
rect 35992 28203 36044 28212
rect 35992 28169 36001 28203
rect 36001 28169 36035 28203
rect 36035 28169 36044 28203
rect 35992 28160 36044 28169
rect 26332 28024 26384 28076
rect 26976 28024 27028 28076
rect 28172 28067 28224 28076
rect 28172 28033 28206 28067
rect 28206 28033 28224 28067
rect 28172 28024 28224 28033
rect 26516 27956 26568 28008
rect 19984 27888 20036 27940
rect 20260 27888 20312 27940
rect 19616 27820 19668 27872
rect 23020 27820 23072 27872
rect 23480 27820 23532 27872
rect 25228 27888 25280 27940
rect 30196 28067 30248 28076
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 31024 28067 31076 28076
rect 31024 28033 31033 28067
rect 31033 28033 31067 28067
rect 31067 28033 31076 28067
rect 31024 28024 31076 28033
rect 31760 28024 31812 28076
rect 30380 27999 30432 28008
rect 30380 27965 30389 27999
rect 30389 27965 30423 27999
rect 30423 27965 30432 27999
rect 30380 27956 30432 27965
rect 31668 27956 31720 28008
rect 36452 28024 36504 28076
rect 31760 27888 31812 27940
rect 24032 27820 24084 27872
rect 26240 27820 26292 27872
rect 31116 27820 31168 27872
rect 31484 27820 31536 27872
rect 36452 27820 36504 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2044 27616 2096 27668
rect 11796 27616 11848 27668
rect 16212 27616 16264 27668
rect 19892 27659 19944 27668
rect 19892 27625 19901 27659
rect 19901 27625 19935 27659
rect 19935 27625 19944 27659
rect 19892 27616 19944 27625
rect 11152 27591 11204 27600
rect 11152 27557 11161 27591
rect 11161 27557 11195 27591
rect 11195 27557 11204 27591
rect 11152 27548 11204 27557
rect 13360 27591 13412 27600
rect 13360 27557 13369 27591
rect 13369 27557 13403 27591
rect 13403 27557 13412 27591
rect 13360 27548 13412 27557
rect 9588 27523 9640 27532
rect 9588 27489 9597 27523
rect 9597 27489 9631 27523
rect 9631 27489 9640 27523
rect 9588 27480 9640 27489
rect 11060 27480 11112 27532
rect 13084 27523 13136 27532
rect 13084 27489 13093 27523
rect 13093 27489 13127 27523
rect 13127 27489 13136 27523
rect 13084 27480 13136 27489
rect 18420 27523 18472 27532
rect 18420 27489 18429 27523
rect 18429 27489 18463 27523
rect 18463 27489 18472 27523
rect 18420 27480 18472 27489
rect 19432 27523 19484 27532
rect 19432 27489 19441 27523
rect 19441 27489 19475 27523
rect 19475 27489 19484 27523
rect 19432 27480 19484 27489
rect 31024 27616 31076 27668
rect 31668 27616 31720 27668
rect 27804 27548 27856 27600
rect 27988 27548 28040 27600
rect 28540 27591 28592 27600
rect 28540 27557 28549 27591
rect 28549 27557 28583 27591
rect 28583 27557 28592 27591
rect 28540 27548 28592 27557
rect 21272 27480 21324 27532
rect 27436 27523 27488 27532
rect 27436 27489 27445 27523
rect 27445 27489 27479 27523
rect 27479 27489 27488 27523
rect 27436 27480 27488 27489
rect 30380 27480 30432 27532
rect 2412 27412 2464 27464
rect 3608 27412 3660 27464
rect 9404 27412 9456 27464
rect 10784 27455 10836 27464
rect 10784 27421 10793 27455
rect 10793 27421 10827 27455
rect 10827 27421 10836 27455
rect 10784 27412 10836 27421
rect 13912 27412 13964 27464
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 15476 27455 15528 27464
rect 15476 27421 15485 27455
rect 15485 27421 15519 27455
rect 15519 27421 15528 27455
rect 15660 27455 15712 27464
rect 15476 27412 15528 27421
rect 15660 27421 15669 27455
rect 15669 27421 15703 27455
rect 15703 27421 15712 27455
rect 15660 27412 15712 27421
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 19616 27455 19668 27464
rect 15752 27412 15804 27421
rect 19616 27421 19625 27455
rect 19625 27421 19659 27455
rect 19659 27421 19668 27455
rect 19616 27412 19668 27421
rect 20260 27412 20312 27464
rect 20996 27412 21048 27464
rect 23020 27455 23072 27464
rect 18144 27387 18196 27396
rect 18144 27353 18162 27387
rect 18162 27353 18196 27387
rect 18144 27344 18196 27353
rect 20904 27344 20956 27396
rect 15660 27276 15712 27328
rect 19432 27276 19484 27328
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 24032 27455 24084 27464
rect 24032 27421 24041 27455
rect 24041 27421 24075 27455
rect 24075 27421 24084 27455
rect 24032 27412 24084 27421
rect 23572 27344 23624 27396
rect 23756 27344 23808 27396
rect 24860 27344 24912 27396
rect 26700 27412 26752 27464
rect 27344 27455 27396 27464
rect 27344 27421 27353 27455
rect 27353 27421 27387 27455
rect 27387 27421 27396 27455
rect 27344 27412 27396 27421
rect 27528 27412 27580 27464
rect 27712 27412 27764 27464
rect 29092 27412 29144 27464
rect 30196 27412 30248 27464
rect 31116 27480 31168 27532
rect 31392 27455 31444 27464
rect 31392 27421 31401 27455
rect 31401 27421 31435 27455
rect 31435 27421 31444 27455
rect 31392 27412 31444 27421
rect 32496 27480 32548 27532
rect 36452 27523 36504 27532
rect 36452 27489 36461 27523
rect 36461 27489 36495 27523
rect 36495 27489 36504 27523
rect 36452 27480 36504 27489
rect 26056 27344 26108 27396
rect 30656 27344 30708 27396
rect 31760 27344 31812 27396
rect 37556 27344 37608 27396
rect 38292 27387 38344 27396
rect 38292 27353 38301 27387
rect 38301 27353 38335 27387
rect 38335 27353 38344 27387
rect 38292 27344 38344 27353
rect 21732 27276 21784 27328
rect 22928 27319 22980 27328
rect 22928 27285 22943 27319
rect 22943 27285 22977 27319
rect 22977 27285 22980 27319
rect 23848 27319 23900 27328
rect 22928 27276 22980 27285
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 24032 27276 24084 27328
rect 25688 27276 25740 27328
rect 26424 27276 26476 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 18144 27072 18196 27124
rect 20260 27072 20312 27124
rect 25688 27115 25740 27124
rect 25688 27081 25697 27115
rect 25697 27081 25731 27115
rect 25731 27081 25740 27115
rect 25688 27072 25740 27081
rect 37556 27115 37608 27124
rect 37556 27081 37565 27115
rect 37565 27081 37599 27115
rect 37599 27081 37608 27115
rect 37556 27072 37608 27081
rect 16856 27004 16908 27056
rect 17408 27047 17460 27056
rect 17408 27013 17417 27047
rect 17417 27013 17451 27047
rect 17451 27013 17460 27047
rect 17408 27004 17460 27013
rect 22744 27004 22796 27056
rect 8576 26979 8628 26988
rect 8576 26945 8585 26979
rect 8585 26945 8619 26979
rect 8619 26945 8628 26979
rect 8576 26936 8628 26945
rect 8944 26936 8996 26988
rect 9220 26979 9272 26988
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 9312 26868 9364 26920
rect 12348 26936 12400 26988
rect 12624 26979 12676 26988
rect 12624 26945 12633 26979
rect 12633 26945 12667 26979
rect 12667 26945 12676 26979
rect 12624 26936 12676 26945
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 13912 26868 13964 26920
rect 12716 26800 12768 26852
rect 3976 26732 4028 26784
rect 9404 26775 9456 26784
rect 9404 26741 9413 26775
rect 9413 26741 9447 26775
rect 9447 26741 9456 26775
rect 9404 26732 9456 26741
rect 10876 26732 10928 26784
rect 11980 26732 12032 26784
rect 12348 26732 12400 26784
rect 17224 26800 17276 26852
rect 19248 26936 19300 26988
rect 23480 26979 23532 26988
rect 23480 26945 23489 26979
rect 23489 26945 23523 26979
rect 23523 26945 23532 26979
rect 23480 26936 23532 26945
rect 23848 27004 23900 27056
rect 31760 27004 31812 27056
rect 24860 26936 24912 26988
rect 24952 26936 25004 26988
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 19340 26911 19392 26920
rect 19340 26877 19349 26911
rect 19349 26877 19383 26911
rect 19383 26877 19392 26911
rect 19340 26868 19392 26877
rect 23940 26868 23992 26920
rect 27344 26936 27396 26988
rect 27620 26936 27672 26988
rect 27528 26868 27580 26920
rect 29276 26868 29328 26920
rect 29736 26936 29788 26988
rect 18328 26800 18380 26852
rect 24860 26800 24912 26852
rect 25504 26843 25556 26852
rect 25504 26809 25513 26843
rect 25513 26809 25547 26843
rect 25547 26809 25556 26843
rect 25504 26800 25556 26809
rect 17316 26732 17368 26784
rect 21364 26732 21416 26784
rect 22928 26732 22980 26784
rect 24308 26732 24360 26784
rect 24676 26732 24728 26784
rect 26332 26775 26384 26784
rect 26332 26741 26341 26775
rect 26341 26741 26375 26775
rect 26375 26741 26384 26775
rect 26332 26732 26384 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8760 26528 8812 26580
rect 9220 26528 9272 26580
rect 9588 26571 9640 26580
rect 9588 26537 9597 26571
rect 9597 26537 9631 26571
rect 9631 26537 9640 26571
rect 9588 26528 9640 26537
rect 10784 26528 10836 26580
rect 12808 26571 12860 26580
rect 4068 26460 4120 26512
rect 3976 26435 4028 26444
rect 3976 26401 3985 26435
rect 3985 26401 4019 26435
rect 4019 26401 4028 26435
rect 3976 26392 4028 26401
rect 9404 26435 9456 26444
rect 9404 26401 9413 26435
rect 9413 26401 9447 26435
rect 9447 26401 9456 26435
rect 9404 26392 9456 26401
rect 4160 26299 4212 26308
rect 4160 26265 4169 26299
rect 4169 26265 4203 26299
rect 4203 26265 4212 26299
rect 4160 26256 4212 26265
rect 8944 26324 8996 26376
rect 9588 26324 9640 26376
rect 12808 26537 12817 26571
rect 12817 26537 12851 26571
rect 12851 26537 12860 26571
rect 12808 26528 12860 26537
rect 17408 26571 17460 26580
rect 17408 26537 17417 26571
rect 17417 26537 17451 26571
rect 17451 26537 17460 26571
rect 17408 26528 17460 26537
rect 22744 26528 22796 26580
rect 23940 26528 23992 26580
rect 25780 26571 25832 26580
rect 10784 26367 10836 26376
rect 10784 26333 10793 26367
rect 10793 26333 10827 26367
rect 10827 26333 10836 26367
rect 10784 26324 10836 26333
rect 10876 26367 10928 26376
rect 10876 26333 10885 26367
rect 10885 26333 10919 26367
rect 10919 26333 10928 26367
rect 11980 26367 12032 26376
rect 10876 26324 10928 26333
rect 11980 26333 11989 26367
rect 11989 26333 12023 26367
rect 12023 26333 12032 26367
rect 11980 26324 12032 26333
rect 12164 26367 12216 26376
rect 12164 26333 12173 26367
rect 12173 26333 12207 26367
rect 12207 26333 12216 26367
rect 12624 26392 12676 26444
rect 14280 26367 14332 26376
rect 12164 26324 12216 26333
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 19156 26460 19208 26512
rect 20628 26460 20680 26512
rect 15936 26435 15988 26444
rect 15936 26401 15945 26435
rect 15945 26401 15979 26435
rect 15979 26401 15988 26435
rect 15936 26392 15988 26401
rect 16120 26392 16172 26444
rect 25780 26537 25789 26571
rect 25789 26537 25823 26571
rect 25823 26537 25832 26571
rect 25780 26528 25832 26537
rect 26792 26571 26844 26580
rect 26792 26537 26801 26571
rect 26801 26537 26835 26571
rect 26835 26537 26844 26571
rect 26792 26528 26844 26537
rect 27436 26528 27488 26580
rect 27804 26571 27856 26580
rect 27804 26537 27813 26571
rect 27813 26537 27847 26571
rect 27847 26537 27856 26571
rect 27804 26528 27856 26537
rect 27988 26571 28040 26580
rect 27988 26537 27997 26571
rect 27997 26537 28031 26571
rect 28031 26537 28040 26571
rect 27988 26528 28040 26537
rect 27620 26460 27672 26512
rect 8576 26256 8628 26308
rect 9128 26256 9180 26308
rect 11060 26299 11112 26308
rect 11060 26265 11069 26299
rect 11069 26265 11103 26299
rect 11103 26265 11112 26299
rect 11060 26256 11112 26265
rect 15844 26367 15896 26376
rect 15844 26333 15853 26367
rect 15853 26333 15887 26367
rect 15887 26333 15896 26367
rect 17592 26367 17644 26376
rect 15844 26324 15896 26333
rect 17592 26333 17601 26367
rect 17601 26333 17635 26367
rect 17635 26333 17644 26367
rect 17592 26324 17644 26333
rect 18604 26324 18656 26376
rect 20260 26324 20312 26376
rect 20904 26324 20956 26376
rect 21824 26324 21876 26376
rect 19984 26256 20036 26308
rect 30288 26528 30340 26580
rect 23572 26324 23624 26376
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 24308 26324 24360 26376
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 27344 26324 27396 26376
rect 27896 26367 27948 26376
rect 27896 26333 27905 26367
rect 27905 26333 27939 26367
rect 27939 26333 27948 26367
rect 27896 26324 27948 26333
rect 28264 26324 28316 26376
rect 28632 26324 28684 26376
rect 29000 26367 29052 26376
rect 29000 26333 29009 26367
rect 29009 26333 29043 26367
rect 29043 26333 29052 26367
rect 29000 26324 29052 26333
rect 33876 26460 33928 26512
rect 24952 26256 25004 26308
rect 26332 26256 26384 26308
rect 29736 26256 29788 26308
rect 33600 26324 33652 26376
rect 12900 26188 12952 26240
rect 15752 26188 15804 26240
rect 17408 26188 17460 26240
rect 19432 26188 19484 26240
rect 26240 26188 26292 26240
rect 27068 26188 27120 26240
rect 29092 26231 29144 26240
rect 29092 26197 29101 26231
rect 29101 26197 29135 26231
rect 29135 26197 29144 26231
rect 29092 26188 29144 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 8852 25984 8904 26036
rect 11060 25984 11112 26036
rect 8760 25959 8812 25968
rect 8760 25925 8769 25959
rect 8769 25925 8803 25959
rect 8803 25925 8812 25959
rect 8760 25916 8812 25925
rect 12716 25984 12768 26036
rect 14280 25984 14332 26036
rect 15936 25984 15988 26036
rect 17224 26027 17276 26036
rect 17224 25993 17233 26027
rect 17233 25993 17267 26027
rect 17267 25993 17276 26027
rect 17224 25984 17276 25993
rect 17592 25959 17644 25968
rect 9312 25848 9364 25900
rect 9588 25891 9640 25900
rect 9588 25857 9597 25891
rect 9597 25857 9631 25891
rect 9631 25857 9640 25891
rect 9588 25848 9640 25857
rect 17592 25925 17601 25959
rect 17601 25925 17635 25959
rect 17635 25925 17644 25959
rect 17592 25916 17644 25925
rect 18052 25916 18104 25968
rect 26332 25984 26384 26036
rect 27528 25984 27580 26036
rect 20628 25959 20680 25968
rect 20628 25925 20646 25959
rect 20646 25925 20680 25959
rect 20628 25916 20680 25925
rect 26240 25916 26292 25968
rect 11796 25848 11848 25900
rect 12440 25891 12492 25900
rect 12440 25857 12449 25891
rect 12449 25857 12483 25891
rect 12483 25857 12492 25891
rect 12440 25848 12492 25857
rect 12716 25891 12768 25900
rect 12716 25857 12750 25891
rect 12750 25857 12768 25891
rect 12716 25848 12768 25857
rect 15844 25848 15896 25900
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 22652 25848 22704 25900
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 27620 25916 27672 25968
rect 29092 25916 29144 25968
rect 15200 25780 15252 25832
rect 16120 25780 16172 25832
rect 26332 25780 26384 25832
rect 26792 25780 26844 25832
rect 27804 25891 27856 25900
rect 27804 25857 27813 25891
rect 27813 25857 27847 25891
rect 27847 25857 27856 25891
rect 27804 25848 27856 25857
rect 28264 25848 28316 25900
rect 30748 25891 30800 25900
rect 27620 25780 27672 25832
rect 28080 25780 28132 25832
rect 30748 25857 30757 25891
rect 30757 25857 30791 25891
rect 30791 25857 30800 25891
rect 30748 25848 30800 25857
rect 38384 25848 38436 25900
rect 14280 25712 14332 25764
rect 14924 25712 14976 25764
rect 18604 25712 18656 25764
rect 21824 25712 21876 25764
rect 25228 25712 25280 25764
rect 17408 25687 17460 25696
rect 17408 25653 17417 25687
rect 17417 25653 17451 25687
rect 17451 25653 17460 25687
rect 17408 25644 17460 25653
rect 19432 25644 19484 25696
rect 19892 25644 19944 25696
rect 26148 25644 26200 25696
rect 26516 25687 26568 25696
rect 26516 25653 26525 25687
rect 26525 25653 26559 25687
rect 26559 25653 26568 25687
rect 26516 25644 26568 25653
rect 26608 25644 26660 25696
rect 31392 25644 31444 25696
rect 38108 25644 38160 25696
rect 38292 25687 38344 25696
rect 38292 25653 38301 25687
rect 38301 25653 38335 25687
rect 38335 25653 38344 25687
rect 38292 25644 38344 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4068 25483 4120 25492
rect 4068 25449 4077 25483
rect 4077 25449 4111 25483
rect 4111 25449 4120 25483
rect 4068 25440 4120 25449
rect 12716 25483 12768 25492
rect 12716 25449 12725 25483
rect 12725 25449 12759 25483
rect 12759 25449 12768 25483
rect 12716 25440 12768 25449
rect 14924 25483 14976 25492
rect 14924 25449 14933 25483
rect 14933 25449 14967 25483
rect 14967 25449 14976 25483
rect 14924 25440 14976 25449
rect 15752 25440 15804 25492
rect 18052 25483 18104 25492
rect 18052 25449 18061 25483
rect 18061 25449 18095 25483
rect 18095 25449 18104 25483
rect 18052 25440 18104 25449
rect 19984 25440 20036 25492
rect 24032 25440 24084 25492
rect 24584 25483 24636 25492
rect 24584 25449 24593 25483
rect 24593 25449 24627 25483
rect 24627 25449 24636 25483
rect 24584 25440 24636 25449
rect 24768 25372 24820 25424
rect 27712 25440 27764 25492
rect 30380 25440 30432 25492
rect 31852 25372 31904 25424
rect 15936 25304 15988 25356
rect 17132 25304 17184 25356
rect 18512 25304 18564 25356
rect 19156 25304 19208 25356
rect 19432 25304 19484 25356
rect 21824 25304 21876 25356
rect 26516 25304 26568 25356
rect 37832 25347 37884 25356
rect 37832 25313 37841 25347
rect 37841 25313 37875 25347
rect 37875 25313 37884 25347
rect 37832 25304 37884 25313
rect 38108 25347 38160 25356
rect 38108 25313 38117 25347
rect 38117 25313 38151 25347
rect 38151 25313 38160 25347
rect 38108 25304 38160 25313
rect 38292 25347 38344 25356
rect 38292 25313 38301 25347
rect 38301 25313 38335 25347
rect 38335 25313 38344 25347
rect 38292 25304 38344 25313
rect 3884 25236 3936 25288
rect 12900 25279 12952 25288
rect 12900 25245 12909 25279
rect 12909 25245 12943 25279
rect 12943 25245 12952 25279
rect 12900 25236 12952 25245
rect 15200 25236 15252 25288
rect 17776 25236 17828 25288
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 18604 25236 18656 25288
rect 17132 25168 17184 25220
rect 18420 25168 18472 25220
rect 19892 25279 19944 25288
rect 19892 25245 19901 25279
rect 19901 25245 19935 25279
rect 19935 25245 19944 25279
rect 19892 25236 19944 25245
rect 20812 25236 20864 25288
rect 22284 25236 22336 25288
rect 24768 25279 24820 25288
rect 24768 25245 24777 25279
rect 24777 25245 24811 25279
rect 24811 25245 24820 25279
rect 24768 25236 24820 25245
rect 26608 25236 26660 25288
rect 27068 25279 27120 25288
rect 27068 25245 27077 25279
rect 27077 25245 27111 25279
rect 27111 25245 27120 25279
rect 27068 25236 27120 25245
rect 16672 25100 16724 25152
rect 21272 25143 21324 25152
rect 21272 25109 21281 25143
rect 21281 25109 21315 25143
rect 21315 25109 21324 25143
rect 21272 25100 21324 25109
rect 22468 25168 22520 25220
rect 22836 25168 22888 25220
rect 26792 25168 26844 25220
rect 27252 25279 27304 25288
rect 27252 25245 27261 25279
rect 27261 25245 27295 25279
rect 27295 25245 27304 25279
rect 27252 25236 27304 25245
rect 29092 25236 29144 25288
rect 31392 25236 31444 25288
rect 31484 25279 31536 25288
rect 31484 25245 31493 25279
rect 31493 25245 31527 25279
rect 31527 25245 31536 25279
rect 31484 25236 31536 25245
rect 23204 25100 23256 25152
rect 30656 25100 30708 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 23204 24896 23256 24948
rect 26332 24939 26384 24948
rect 9404 24871 9456 24880
rect 9404 24837 9413 24871
rect 9413 24837 9447 24871
rect 9447 24837 9456 24871
rect 9404 24828 9456 24837
rect 9772 24828 9824 24880
rect 23664 24828 23716 24880
rect 24860 24871 24912 24880
rect 26332 24905 26341 24939
rect 26341 24905 26375 24939
rect 26375 24905 26384 24939
rect 26332 24896 26384 24905
rect 30564 24896 30616 24948
rect 31484 24896 31536 24948
rect 24860 24837 24885 24871
rect 24885 24837 24912 24871
rect 24860 24828 24912 24837
rect 4068 24735 4120 24744
rect 4068 24701 4077 24735
rect 4077 24701 4111 24735
rect 4111 24701 4120 24735
rect 4068 24692 4120 24701
rect 5448 24735 5500 24744
rect 5448 24701 5457 24735
rect 5457 24701 5491 24735
rect 5491 24701 5500 24735
rect 5448 24692 5500 24701
rect 4804 24624 4856 24676
rect 16028 24803 16080 24812
rect 16028 24769 16037 24803
rect 16037 24769 16071 24803
rect 16071 24769 16080 24803
rect 16028 24760 16080 24769
rect 13728 24692 13780 24744
rect 14372 24735 14424 24744
rect 14372 24701 14381 24735
rect 14381 24701 14415 24735
rect 14415 24701 14424 24735
rect 14372 24692 14424 24701
rect 8576 24556 8628 24608
rect 10416 24599 10468 24608
rect 10416 24565 10425 24599
rect 10425 24565 10459 24599
rect 10459 24565 10468 24599
rect 10416 24556 10468 24565
rect 17500 24556 17552 24608
rect 17960 24760 18012 24812
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 22836 24803 22888 24812
rect 22836 24769 22845 24803
rect 22845 24769 22879 24803
rect 22879 24769 22888 24803
rect 22836 24760 22888 24769
rect 26516 24760 26568 24812
rect 26700 24828 26752 24880
rect 27252 24828 27304 24880
rect 27344 24803 27396 24812
rect 27344 24769 27353 24803
rect 27353 24769 27387 24803
rect 27387 24769 27396 24803
rect 27344 24760 27396 24769
rect 27988 24760 28040 24812
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 28908 24760 28960 24812
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 29736 24760 29788 24812
rect 22284 24692 22336 24744
rect 26792 24692 26844 24744
rect 27620 24735 27672 24744
rect 27620 24701 27629 24735
rect 27629 24701 27663 24735
rect 27663 24701 27672 24735
rect 27620 24692 27672 24701
rect 28172 24735 28224 24744
rect 28172 24701 28181 24735
rect 28181 24701 28215 24735
rect 28215 24701 28224 24735
rect 28172 24692 28224 24701
rect 30656 24760 30708 24812
rect 31116 24803 31168 24812
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 31392 24803 31444 24812
rect 31392 24769 31401 24803
rect 31401 24769 31435 24803
rect 31435 24769 31444 24803
rect 31392 24760 31444 24769
rect 37280 24760 37332 24812
rect 20352 24624 20404 24676
rect 30196 24692 30248 24744
rect 29000 24624 29052 24676
rect 21364 24599 21416 24608
rect 21364 24565 21373 24599
rect 21373 24565 21407 24599
rect 21407 24565 21416 24599
rect 21364 24556 21416 24565
rect 24768 24556 24820 24608
rect 25136 24556 25188 24608
rect 25504 24599 25556 24608
rect 25504 24565 25513 24599
rect 25513 24565 25547 24599
rect 25547 24565 25556 24599
rect 25504 24556 25556 24565
rect 26332 24556 26384 24608
rect 26884 24556 26936 24608
rect 28632 24556 28684 24608
rect 38108 24556 38160 24608
rect 38292 24599 38344 24608
rect 38292 24565 38301 24599
rect 38301 24565 38335 24599
rect 38335 24565 38344 24599
rect 38292 24556 38344 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4068 24395 4120 24404
rect 4068 24361 4077 24395
rect 4077 24361 4111 24395
rect 4111 24361 4120 24395
rect 4068 24352 4120 24361
rect 9404 24352 9456 24404
rect 11796 24352 11848 24404
rect 13728 24395 13780 24404
rect 13728 24361 13737 24395
rect 13737 24361 13771 24395
rect 13771 24361 13780 24395
rect 13728 24352 13780 24361
rect 14280 24352 14332 24404
rect 19340 24352 19392 24404
rect 22468 24395 22520 24404
rect 22468 24361 22477 24395
rect 22477 24361 22511 24395
rect 22511 24361 22520 24395
rect 22468 24352 22520 24361
rect 25504 24352 25556 24404
rect 26516 24395 26568 24404
rect 26516 24361 26525 24395
rect 26525 24361 26559 24395
rect 26559 24361 26568 24395
rect 26516 24352 26568 24361
rect 26700 24395 26752 24404
rect 26700 24361 26709 24395
rect 26709 24361 26743 24395
rect 26743 24361 26752 24395
rect 26700 24352 26752 24361
rect 28908 24395 28960 24404
rect 28908 24361 28917 24395
rect 28917 24361 28951 24395
rect 28951 24361 28960 24395
rect 28908 24352 28960 24361
rect 29736 24395 29788 24404
rect 29736 24361 29745 24395
rect 29745 24361 29779 24395
rect 29779 24361 29788 24395
rect 29736 24352 29788 24361
rect 12532 24216 12584 24268
rect 3884 24148 3936 24200
rect 8576 24191 8628 24200
rect 8576 24157 8585 24191
rect 8585 24157 8619 24191
rect 8619 24157 8628 24191
rect 8576 24148 8628 24157
rect 10232 24148 10284 24200
rect 12348 24148 12400 24200
rect 14096 24148 14148 24200
rect 10048 24080 10100 24132
rect 10416 24080 10468 24132
rect 10692 24080 10744 24132
rect 16672 24123 16724 24132
rect 9036 24012 9088 24064
rect 9128 24012 9180 24064
rect 13360 24012 13412 24064
rect 15200 24012 15252 24064
rect 16120 24055 16172 24064
rect 16120 24021 16129 24055
rect 16129 24021 16163 24055
rect 16163 24021 16172 24055
rect 16120 24012 16172 24021
rect 16672 24089 16681 24123
rect 16681 24089 16715 24123
rect 16715 24089 16724 24123
rect 16672 24080 16724 24089
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 16948 24012 17000 24064
rect 17592 24080 17644 24132
rect 18512 24148 18564 24200
rect 18788 24191 18840 24200
rect 18788 24157 18797 24191
rect 18797 24157 18831 24191
rect 18831 24157 18840 24191
rect 18788 24148 18840 24157
rect 20076 24148 20128 24200
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 20812 24012 20864 24064
rect 22652 24216 22704 24268
rect 28080 24284 28132 24336
rect 25136 24259 25188 24268
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23204 24080 23256 24132
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 25136 24225 25145 24259
rect 25145 24225 25179 24259
rect 25179 24225 25188 24259
rect 25136 24216 25188 24225
rect 26792 24259 26844 24268
rect 26792 24225 26801 24259
rect 26801 24225 26835 24259
rect 26835 24225 26844 24259
rect 26792 24216 26844 24225
rect 28632 24259 28684 24268
rect 28632 24225 28641 24259
rect 28641 24225 28675 24259
rect 28675 24225 28684 24259
rect 28632 24216 28684 24225
rect 23756 24148 23808 24157
rect 26884 24191 26936 24200
rect 26884 24157 26893 24191
rect 26893 24157 26927 24191
rect 26927 24157 26936 24191
rect 26884 24148 26936 24157
rect 27344 24148 27396 24200
rect 27988 24148 28040 24200
rect 28264 24148 28316 24200
rect 29184 24148 29236 24200
rect 30656 24216 30708 24268
rect 37832 24259 37884 24268
rect 37832 24225 37841 24259
rect 37841 24225 37875 24259
rect 37875 24225 37884 24259
rect 37832 24216 37884 24225
rect 38108 24259 38160 24268
rect 38108 24225 38117 24259
rect 38117 24225 38151 24259
rect 38151 24225 38160 24259
rect 38108 24216 38160 24225
rect 38292 24259 38344 24268
rect 38292 24225 38301 24259
rect 38301 24225 38335 24259
rect 38335 24225 38344 24259
rect 38292 24216 38344 24225
rect 30196 24191 30248 24200
rect 30196 24157 30205 24191
rect 30205 24157 30239 24191
rect 30239 24157 30248 24191
rect 30196 24148 30248 24157
rect 23572 24012 23624 24064
rect 24768 24012 24820 24064
rect 24860 24012 24912 24064
rect 31116 24080 31168 24132
rect 30288 24012 30340 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3884 23808 3936 23860
rect 13820 23808 13872 23860
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 10048 23783 10100 23792
rect 10048 23749 10075 23783
rect 10075 23749 10100 23783
rect 10048 23740 10100 23749
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 9128 23672 9180 23724
rect 9772 23672 9824 23724
rect 10140 23672 10192 23724
rect 11796 23740 11848 23792
rect 12256 23783 12308 23792
rect 12256 23749 12265 23783
rect 12265 23749 12299 23783
rect 12299 23749 12308 23783
rect 12256 23740 12308 23749
rect 16948 23808 17000 23860
rect 17592 23808 17644 23860
rect 18788 23808 18840 23860
rect 20720 23808 20772 23860
rect 23940 23808 23992 23860
rect 29184 23851 29236 23860
rect 29184 23817 29193 23851
rect 29193 23817 29227 23851
rect 29227 23817 29236 23851
rect 29184 23808 29236 23817
rect 12348 23672 12400 23724
rect 15476 23740 15528 23792
rect 18144 23740 18196 23792
rect 20904 23783 20956 23792
rect 20904 23749 20913 23783
rect 20913 23749 20947 23783
rect 20947 23749 20956 23783
rect 20904 23740 20956 23749
rect 22284 23740 22336 23792
rect 24952 23740 25004 23792
rect 27804 23740 27856 23792
rect 29092 23740 29144 23792
rect 29736 23740 29788 23792
rect 35716 23783 35768 23792
rect 35716 23749 35725 23783
rect 35725 23749 35759 23783
rect 35759 23749 35768 23783
rect 35716 23740 35768 23749
rect 13360 23715 13412 23724
rect 13360 23681 13369 23715
rect 13369 23681 13403 23715
rect 13403 23681 13412 23715
rect 14280 23715 14332 23724
rect 13360 23672 13412 23681
rect 14280 23681 14289 23715
rect 14289 23681 14323 23715
rect 14323 23681 14332 23715
rect 14280 23672 14332 23681
rect 13912 23604 13964 23656
rect 14188 23604 14240 23656
rect 15660 23672 15712 23724
rect 18420 23672 18472 23724
rect 22100 23715 22152 23724
rect 22100 23681 22109 23715
rect 22109 23681 22143 23715
rect 22143 23681 22152 23715
rect 22100 23672 22152 23681
rect 24768 23715 24820 23724
rect 24768 23681 24802 23715
rect 24802 23681 24820 23715
rect 24768 23672 24820 23681
rect 26976 23672 27028 23724
rect 18144 23604 18196 23656
rect 10876 23536 10928 23588
rect 8852 23468 8904 23520
rect 10324 23468 10376 23520
rect 13452 23511 13504 23520
rect 13452 23477 13461 23511
rect 13461 23477 13495 23511
rect 13495 23477 13504 23511
rect 13452 23468 13504 23477
rect 17684 23536 17736 23588
rect 20628 23579 20680 23588
rect 20628 23545 20637 23579
rect 20637 23545 20671 23579
rect 20671 23545 20680 23579
rect 20628 23536 20680 23545
rect 22192 23604 22244 23656
rect 27988 23604 28040 23656
rect 33876 23715 33928 23724
rect 33876 23681 33885 23715
rect 33885 23681 33919 23715
rect 33919 23681 33928 23715
rect 33876 23672 33928 23681
rect 34060 23647 34112 23656
rect 34060 23613 34069 23647
rect 34069 23613 34103 23647
rect 34103 23613 34112 23647
rect 34060 23604 34112 23613
rect 16488 23468 16540 23520
rect 22836 23468 22888 23520
rect 30656 23536 30708 23588
rect 30932 23536 30984 23588
rect 26332 23468 26384 23520
rect 27896 23468 27948 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 10140 23307 10192 23316
rect 10140 23273 10149 23307
rect 10149 23273 10183 23307
rect 10183 23273 10192 23307
rect 10140 23264 10192 23273
rect 14372 23307 14424 23316
rect 14372 23273 14381 23307
rect 14381 23273 14415 23307
rect 14415 23273 14424 23307
rect 14372 23264 14424 23273
rect 15844 23264 15896 23316
rect 16488 23264 16540 23316
rect 20076 23264 20128 23316
rect 34060 23264 34112 23316
rect 13728 23196 13780 23248
rect 14280 23196 14332 23248
rect 2412 23060 2464 23112
rect 2596 23060 2648 23112
rect 3700 23060 3752 23112
rect 9036 23060 9088 23112
rect 9588 23103 9640 23112
rect 9588 23069 9597 23103
rect 9597 23069 9631 23103
rect 9631 23069 9640 23103
rect 9588 23060 9640 23069
rect 10324 23128 10376 23180
rect 10140 23060 10192 23112
rect 10692 23060 10744 23112
rect 10876 23060 10928 23112
rect 17132 23128 17184 23180
rect 12256 23060 12308 23112
rect 3516 22924 3568 22976
rect 10048 22924 10100 22976
rect 12348 22992 12400 23044
rect 13820 23060 13872 23112
rect 16120 23060 16172 23112
rect 18420 23196 18472 23248
rect 20168 23239 20220 23248
rect 20168 23205 20177 23239
rect 20177 23205 20211 23239
rect 20211 23205 20220 23239
rect 20168 23196 20220 23205
rect 22100 23196 22152 23248
rect 26792 23239 26844 23248
rect 26792 23205 26801 23239
rect 26801 23205 26835 23239
rect 26835 23205 26844 23239
rect 26792 23196 26844 23205
rect 21088 23128 21140 23180
rect 17776 23103 17828 23112
rect 17776 23069 17785 23103
rect 17785 23069 17819 23103
rect 17819 23069 17828 23103
rect 17776 23060 17828 23069
rect 18052 23060 18104 23112
rect 17868 22992 17920 23044
rect 14740 22924 14792 22976
rect 17040 22967 17092 22976
rect 17040 22933 17065 22967
rect 17065 22933 17092 22967
rect 17040 22924 17092 22933
rect 17684 22924 17736 22976
rect 20352 22992 20404 23044
rect 22284 23128 22336 23180
rect 23572 23128 23624 23180
rect 24860 23128 24912 23180
rect 26332 23171 26384 23180
rect 26332 23137 26341 23171
rect 26341 23137 26375 23171
rect 26375 23137 26384 23171
rect 26332 23128 26384 23137
rect 30380 23128 30432 23180
rect 23664 23103 23716 23112
rect 23664 23069 23673 23103
rect 23673 23069 23707 23103
rect 23707 23069 23716 23103
rect 23664 23060 23716 23069
rect 24308 23060 24360 23112
rect 26976 23060 27028 23112
rect 30748 23060 30800 23112
rect 31852 23103 31904 23112
rect 31852 23069 31861 23103
rect 31861 23069 31895 23103
rect 31895 23069 31904 23103
rect 31852 23060 31904 23069
rect 33876 23060 33928 23112
rect 38292 23060 38344 23112
rect 24216 22992 24268 23044
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 21916 22924 21968 22976
rect 22744 22967 22796 22976
rect 22744 22933 22753 22967
rect 22753 22933 22787 22967
rect 22787 22933 22796 22967
rect 22744 22924 22796 22933
rect 23756 22924 23808 22976
rect 31024 22924 31076 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3516 22695 3568 22704
rect 3516 22661 3525 22695
rect 3525 22661 3559 22695
rect 3559 22661 3568 22695
rect 3516 22652 3568 22661
rect 3700 22627 3752 22636
rect 3700 22593 3709 22627
rect 3709 22593 3743 22627
rect 3743 22593 3752 22627
rect 13728 22720 13780 22772
rect 15476 22763 15528 22772
rect 15476 22729 15485 22763
rect 15485 22729 15519 22763
rect 15519 22729 15528 22763
rect 15476 22720 15528 22729
rect 17776 22720 17828 22772
rect 18236 22763 18288 22772
rect 18236 22729 18245 22763
rect 18245 22729 18279 22763
rect 18279 22729 18288 22763
rect 18236 22720 18288 22729
rect 3700 22584 3752 22593
rect 12440 22584 12492 22636
rect 13452 22584 13504 22636
rect 14832 22584 14884 22636
rect 1860 22559 1912 22568
rect 1860 22525 1869 22559
rect 1869 22525 1903 22559
rect 1903 22525 1912 22559
rect 1860 22516 1912 22525
rect 9588 22516 9640 22568
rect 12716 22516 12768 22568
rect 15660 22584 15712 22636
rect 16120 22652 16172 22704
rect 17592 22652 17644 22704
rect 17868 22652 17920 22704
rect 21916 22720 21968 22772
rect 30564 22763 30616 22772
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 17408 22584 17460 22636
rect 9864 22448 9916 22500
rect 22284 22652 22336 22704
rect 22744 22652 22796 22704
rect 19984 22516 20036 22568
rect 20536 22627 20588 22636
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 22192 22627 22244 22636
rect 20720 22584 20772 22593
rect 21364 22516 21416 22568
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 30564 22729 30573 22763
rect 30573 22729 30607 22763
rect 30607 22729 30616 22763
rect 30564 22720 30616 22729
rect 24768 22695 24820 22704
rect 24768 22661 24777 22695
rect 24777 22661 24811 22695
rect 24811 22661 24820 22695
rect 24768 22652 24820 22661
rect 29552 22584 29604 22636
rect 30380 22584 30432 22636
rect 31024 22627 31076 22636
rect 31024 22593 31033 22627
rect 31033 22593 31067 22627
rect 31067 22593 31076 22627
rect 31024 22584 31076 22593
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 37740 22584 37792 22636
rect 29276 22516 29328 22568
rect 30656 22516 30708 22568
rect 23572 22491 23624 22500
rect 23572 22457 23581 22491
rect 23581 22457 23615 22491
rect 23615 22457 23624 22491
rect 23572 22448 23624 22457
rect 24768 22448 24820 22500
rect 25872 22448 25924 22500
rect 15844 22380 15896 22432
rect 18420 22380 18472 22432
rect 23388 22380 23440 22432
rect 30380 22423 30432 22432
rect 30380 22389 30389 22423
rect 30389 22389 30423 22423
rect 30423 22389 30432 22423
rect 30380 22380 30432 22389
rect 38108 22380 38160 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 13084 22176 13136 22228
rect 14096 22176 14148 22228
rect 15016 22176 15068 22228
rect 15476 22176 15528 22228
rect 20536 22176 20588 22228
rect 20720 22176 20772 22228
rect 21180 22176 21232 22228
rect 26056 22176 26108 22228
rect 28632 22176 28684 22228
rect 30472 22176 30524 22228
rect 2780 22083 2832 22092
rect 2780 22049 2789 22083
rect 2789 22049 2823 22083
rect 2823 22049 2832 22083
rect 2780 22040 2832 22049
rect 8668 22040 8720 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 14188 22040 14240 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 15660 22083 15712 22092
rect 14740 22040 14792 22049
rect 15660 22049 15669 22083
rect 15669 22049 15703 22083
rect 15703 22049 15712 22083
rect 15660 22040 15712 22049
rect 17408 22083 17460 22092
rect 17408 22049 17417 22083
rect 17417 22049 17451 22083
rect 17451 22049 17460 22083
rect 17408 22040 17460 22049
rect 17868 22083 17920 22092
rect 17868 22049 17877 22083
rect 17877 22049 17911 22083
rect 17911 22049 17920 22083
rect 17868 22040 17920 22049
rect 24216 22040 24268 22092
rect 12716 21972 12768 22024
rect 13176 21972 13228 22024
rect 13452 22015 13504 22024
rect 13452 21981 13461 22015
rect 13461 21981 13495 22015
rect 13495 21981 13504 22015
rect 14924 22015 14976 22024
rect 13452 21972 13504 21981
rect 14924 21981 14933 22015
rect 14933 21981 14967 22015
rect 14967 21981 14976 22015
rect 14924 21972 14976 21981
rect 15016 21972 15068 22024
rect 20076 22015 20128 22024
rect 2412 21904 2464 21956
rect 10048 21904 10100 21956
rect 12992 21904 13044 21956
rect 14372 21904 14424 21956
rect 15568 21947 15620 21956
rect 15568 21913 15577 21947
rect 15577 21913 15611 21947
rect 15611 21913 15620 21947
rect 15568 21904 15620 21913
rect 12440 21836 12492 21888
rect 15108 21879 15160 21888
rect 15108 21845 15117 21879
rect 15117 21845 15151 21879
rect 15151 21845 15160 21879
rect 15108 21836 15160 21845
rect 20076 21981 20085 22015
rect 20085 21981 20119 22015
rect 20119 21981 20128 22015
rect 20076 21972 20128 21981
rect 20904 21972 20956 22024
rect 21272 21972 21324 22024
rect 23756 21972 23808 22024
rect 24860 22015 24912 22024
rect 18512 21904 18564 21956
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 24860 21972 24912 21981
rect 25872 22040 25924 22092
rect 27344 22083 27396 22092
rect 27344 22049 27353 22083
rect 27353 22049 27387 22083
rect 27387 22049 27396 22083
rect 27344 22040 27396 22049
rect 24124 21904 24176 21956
rect 24400 21904 24452 21956
rect 17500 21836 17552 21888
rect 23664 21836 23716 21888
rect 23940 21836 23992 21888
rect 26240 21879 26292 21888
rect 26240 21845 26249 21879
rect 26249 21845 26283 21879
rect 26283 21845 26292 21879
rect 26240 21836 26292 21845
rect 27160 22015 27212 22024
rect 27160 21981 27169 22015
rect 27169 21981 27203 22015
rect 27203 21981 27212 22015
rect 27160 21972 27212 21981
rect 37188 22083 37240 22092
rect 37188 22049 37197 22083
rect 37197 22049 37231 22083
rect 37231 22049 37240 22083
rect 37188 22040 37240 22049
rect 38108 22083 38160 22092
rect 38108 22049 38117 22083
rect 38117 22049 38151 22083
rect 38151 22049 38160 22083
rect 38108 22040 38160 22049
rect 38292 22083 38344 22092
rect 38292 22049 38301 22083
rect 38301 22049 38335 22083
rect 38335 22049 38344 22083
rect 38292 22040 38344 22049
rect 27712 21972 27764 22024
rect 29644 21904 29696 21956
rect 27804 21836 27856 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2412 21675 2464 21684
rect 2412 21641 2421 21675
rect 2421 21641 2455 21675
rect 2455 21641 2464 21675
rect 2412 21632 2464 21641
rect 1584 21496 1636 21548
rect 2688 21496 2740 21548
rect 2780 21496 2832 21548
rect 8668 21496 8720 21548
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 9128 21496 9180 21548
rect 12440 21564 12492 21616
rect 15568 21632 15620 21684
rect 17224 21564 17276 21616
rect 11980 21496 12032 21548
rect 13820 21496 13872 21548
rect 14096 21539 14148 21548
rect 14096 21505 14105 21539
rect 14105 21505 14139 21539
rect 14139 21505 14148 21539
rect 14096 21496 14148 21505
rect 14372 21496 14424 21548
rect 15108 21496 15160 21548
rect 15936 21496 15988 21548
rect 17960 21564 18012 21616
rect 3608 21428 3660 21480
rect 9588 21428 9640 21480
rect 12992 21471 13044 21480
rect 12992 21437 13001 21471
rect 13001 21437 13035 21471
rect 13035 21437 13044 21471
rect 12992 21428 13044 21437
rect 14464 21428 14516 21480
rect 14924 21428 14976 21480
rect 15476 21428 15528 21480
rect 13820 21360 13872 21412
rect 14188 21360 14240 21412
rect 15200 21360 15252 21412
rect 19800 21496 19852 21548
rect 20904 21632 20956 21684
rect 21364 21675 21416 21684
rect 21364 21641 21373 21675
rect 21373 21641 21407 21675
rect 21407 21641 21416 21675
rect 21364 21632 21416 21641
rect 24032 21632 24084 21684
rect 24400 21675 24452 21684
rect 23204 21564 23256 21616
rect 24400 21641 24409 21675
rect 24409 21641 24443 21675
rect 24443 21641 24452 21675
rect 24400 21632 24452 21641
rect 24860 21632 24912 21684
rect 27712 21632 27764 21684
rect 29644 21675 29696 21684
rect 29644 21641 29653 21675
rect 29653 21641 29687 21675
rect 29687 21641 29696 21675
rect 29644 21632 29696 21641
rect 20352 21496 20404 21548
rect 22652 21539 22704 21548
rect 3240 21292 3292 21344
rect 9680 21335 9732 21344
rect 9680 21301 9689 21335
rect 9689 21301 9723 21335
rect 9723 21301 9732 21335
rect 9680 21292 9732 21301
rect 12348 21292 12400 21344
rect 13176 21335 13228 21344
rect 13176 21301 13185 21335
rect 13185 21301 13219 21335
rect 13219 21301 13228 21335
rect 13176 21292 13228 21301
rect 13268 21292 13320 21344
rect 15844 21292 15896 21344
rect 17132 21292 17184 21344
rect 17776 21360 17828 21412
rect 20260 21360 20312 21412
rect 21916 21360 21968 21412
rect 18236 21292 18288 21344
rect 18788 21292 18840 21344
rect 19340 21292 19392 21344
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 23756 21539 23808 21548
rect 23756 21505 23765 21539
rect 23765 21505 23799 21539
rect 23799 21505 23808 21539
rect 23756 21496 23808 21505
rect 23940 21539 23992 21548
rect 23940 21505 23949 21539
rect 23949 21505 23983 21539
rect 23983 21505 23992 21539
rect 23940 21496 23992 21505
rect 27160 21564 27212 21616
rect 35440 21607 35492 21616
rect 35440 21573 35449 21607
rect 35449 21573 35483 21607
rect 35483 21573 35492 21607
rect 35440 21564 35492 21573
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 26700 21496 26752 21548
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 27988 21539 28040 21548
rect 27988 21505 28022 21539
rect 28022 21505 28040 21539
rect 27988 21496 28040 21505
rect 29552 21539 29604 21548
rect 29552 21505 29561 21539
rect 29561 21505 29595 21539
rect 29595 21505 29604 21539
rect 29552 21496 29604 21505
rect 30380 21496 30432 21548
rect 32956 21539 33008 21548
rect 32956 21505 32965 21539
rect 32965 21505 32999 21539
rect 32999 21505 33008 21539
rect 32956 21496 33008 21505
rect 33600 21539 33652 21548
rect 33600 21505 33609 21539
rect 33609 21505 33643 21539
rect 33643 21505 33652 21539
rect 33600 21496 33652 21505
rect 23572 21428 23624 21480
rect 23664 21360 23716 21412
rect 27436 21292 27488 21344
rect 28448 21292 28500 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9128 21131 9180 21140
rect 9128 21097 9137 21131
rect 9137 21097 9171 21131
rect 9171 21097 9180 21131
rect 9128 21088 9180 21097
rect 13176 21088 13228 21140
rect 17408 21088 17460 21140
rect 20076 21020 20128 21072
rect 22100 21020 22152 21072
rect 1584 20995 1636 21004
rect 1584 20961 1593 20995
rect 1593 20961 1627 20995
rect 1627 20961 1636 20995
rect 1584 20952 1636 20961
rect 3240 20995 3292 21004
rect 3240 20961 3249 20995
rect 3249 20961 3283 20995
rect 3283 20961 3292 20995
rect 3240 20952 3292 20961
rect 8300 20927 8352 20936
rect 3056 20816 3108 20868
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 8668 20952 8720 21004
rect 13452 20952 13504 21004
rect 14648 20995 14700 21004
rect 14648 20961 14657 20995
rect 14657 20961 14691 20995
rect 14691 20961 14700 20995
rect 14648 20952 14700 20961
rect 18788 20952 18840 21004
rect 24860 21088 24912 21140
rect 27988 21131 28040 21140
rect 27988 21097 27997 21131
rect 27997 21097 28031 21131
rect 28031 21097 28040 21131
rect 27988 21088 28040 21097
rect 26240 20952 26292 21004
rect 26700 20995 26752 21004
rect 26700 20961 26709 20995
rect 26709 20961 26743 20995
rect 26743 20961 26752 20995
rect 26700 20952 26752 20961
rect 8852 20884 8904 20936
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 14372 20927 14424 20936
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 14372 20884 14424 20893
rect 14464 20927 14516 20936
rect 14464 20893 14473 20927
rect 14473 20893 14507 20927
rect 14507 20893 14516 20927
rect 17224 20927 17276 20936
rect 14464 20884 14516 20893
rect 17224 20893 17233 20927
rect 17233 20893 17267 20927
rect 17267 20893 17276 20927
rect 17224 20884 17276 20893
rect 17592 20884 17644 20936
rect 18512 20927 18564 20936
rect 9588 20816 9640 20868
rect 9680 20816 9732 20868
rect 10692 20816 10744 20868
rect 12440 20859 12492 20868
rect 12440 20825 12474 20859
rect 12474 20825 12492 20859
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 19984 20884 20036 20936
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 22100 20884 22152 20936
rect 23388 20884 23440 20936
rect 27712 20927 27764 20936
rect 27712 20893 27721 20927
rect 27721 20893 27755 20927
rect 27755 20893 27764 20927
rect 27712 20884 27764 20893
rect 28448 20927 28500 20936
rect 12440 20816 12492 20825
rect 19800 20859 19852 20868
rect 19800 20825 19809 20859
rect 19809 20825 19843 20859
rect 19843 20825 19852 20859
rect 19800 20816 19852 20825
rect 26608 20816 26660 20868
rect 28448 20893 28457 20927
rect 28457 20893 28491 20927
rect 28491 20893 28500 20927
rect 28448 20884 28500 20893
rect 28632 20927 28684 20936
rect 28632 20893 28641 20927
rect 28641 20893 28675 20927
rect 28675 20893 28684 20927
rect 28632 20884 28684 20893
rect 27896 20816 27948 20868
rect 28172 20816 28224 20868
rect 8576 20791 8628 20800
rect 8576 20757 8585 20791
rect 8585 20757 8619 20791
rect 8619 20757 8628 20791
rect 8576 20748 8628 20757
rect 12992 20748 13044 20800
rect 16764 20748 16816 20800
rect 17040 20748 17092 20800
rect 17960 20791 18012 20800
rect 17960 20757 17969 20791
rect 17969 20757 18003 20791
rect 18003 20757 18012 20791
rect 17960 20748 18012 20757
rect 18972 20748 19024 20800
rect 19432 20791 19484 20800
rect 19432 20757 19441 20791
rect 19441 20757 19475 20791
rect 19475 20757 19484 20791
rect 19432 20748 19484 20757
rect 26332 20748 26384 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 8852 20544 8904 20596
rect 12440 20544 12492 20596
rect 16764 20544 16816 20596
rect 16948 20587 17000 20596
rect 16948 20553 16957 20587
rect 16957 20553 16991 20587
rect 16991 20553 17000 20587
rect 16948 20544 17000 20553
rect 17408 20544 17460 20596
rect 20812 20544 20864 20596
rect 1952 20519 2004 20528
rect 1952 20485 1961 20519
rect 1961 20485 1995 20519
rect 1995 20485 2004 20519
rect 1952 20476 2004 20485
rect 8300 20476 8352 20528
rect 8576 20408 8628 20460
rect 2688 20340 2740 20392
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 9128 20315 9180 20324
rect 9128 20281 9137 20315
rect 9137 20281 9171 20315
rect 9171 20281 9180 20315
rect 9128 20272 9180 20281
rect 13176 20476 13228 20528
rect 17960 20476 18012 20528
rect 19432 20476 19484 20528
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 13912 20408 13964 20460
rect 17592 20408 17644 20460
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 18972 20408 19024 20417
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 21180 20451 21232 20460
rect 21180 20417 21198 20451
rect 21198 20417 21232 20451
rect 21180 20408 21232 20417
rect 22008 20408 22060 20460
rect 22284 20451 22336 20460
rect 22284 20417 22293 20451
rect 22293 20417 22327 20451
rect 22327 20417 22336 20451
rect 22284 20408 22336 20417
rect 26240 20408 26292 20460
rect 30564 20587 30616 20596
rect 26700 20476 26752 20528
rect 26516 20408 26568 20460
rect 28080 20408 28132 20460
rect 30564 20553 30573 20587
rect 30573 20553 30607 20587
rect 30607 20553 30616 20587
rect 30564 20544 30616 20553
rect 30932 20544 30984 20596
rect 19984 20340 20036 20392
rect 24032 20340 24084 20392
rect 17960 20272 18012 20324
rect 8668 20204 8720 20256
rect 13084 20204 13136 20256
rect 14648 20204 14700 20256
rect 14832 20204 14884 20256
rect 17132 20204 17184 20256
rect 17316 20204 17368 20256
rect 23204 20272 23256 20324
rect 27896 20340 27948 20392
rect 30472 20451 30524 20460
rect 30472 20417 30514 20451
rect 30514 20417 30524 20451
rect 30472 20408 30524 20417
rect 31116 20408 31168 20460
rect 31668 20340 31720 20392
rect 20720 20204 20772 20256
rect 26976 20204 27028 20256
rect 30840 20272 30892 20324
rect 31576 20315 31628 20324
rect 31576 20281 31585 20315
rect 31585 20281 31619 20315
rect 31619 20281 31628 20315
rect 31576 20272 31628 20281
rect 27988 20247 28040 20256
rect 27988 20213 27997 20247
rect 27997 20213 28031 20247
rect 28031 20213 28040 20247
rect 27988 20204 28040 20213
rect 29920 20204 29972 20256
rect 30564 20204 30616 20256
rect 30748 20204 30800 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2688 20043 2740 20052
rect 2688 20009 2697 20043
rect 2697 20009 2731 20043
rect 2731 20009 2740 20043
rect 2688 20000 2740 20009
rect 3792 20000 3844 20052
rect 3056 19932 3108 19984
rect 4068 19796 4120 19848
rect 5632 19796 5684 19848
rect 11980 19796 12032 19848
rect 14464 19796 14516 19848
rect 4712 19728 4764 19780
rect 16304 20000 16356 20052
rect 18144 20000 18196 20052
rect 16856 19932 16908 19984
rect 21180 20000 21232 20052
rect 26516 20000 26568 20052
rect 27988 20000 28040 20052
rect 31116 20043 31168 20052
rect 31116 20009 31125 20043
rect 31125 20009 31159 20043
rect 31159 20009 31168 20043
rect 31116 20000 31168 20009
rect 31668 20043 31720 20052
rect 31668 20009 31677 20043
rect 31677 20009 31711 20043
rect 31711 20009 31720 20043
rect 31668 20000 31720 20009
rect 16396 19864 16448 19916
rect 17126 19907 17178 19916
rect 17126 19873 17135 19907
rect 17135 19873 17169 19907
rect 17169 19873 17178 19907
rect 17126 19864 17178 19873
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 10232 19660 10284 19712
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 20720 19796 20772 19848
rect 20996 19796 21048 19848
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 27712 19932 27764 19984
rect 27896 19975 27948 19984
rect 27896 19941 27905 19975
rect 27905 19941 27939 19975
rect 27939 19941 27948 19975
rect 27896 19932 27948 19941
rect 23664 19839 23716 19848
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 24032 19839 24084 19848
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 26608 19864 26660 19916
rect 26332 19796 26384 19848
rect 26976 19839 27028 19848
rect 26976 19805 26985 19839
rect 26985 19805 27019 19839
rect 27019 19805 27028 19839
rect 26976 19796 27028 19805
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 27528 19796 27580 19848
rect 27620 19796 27672 19848
rect 30104 19864 30156 19916
rect 31852 19907 31904 19916
rect 31852 19873 31861 19907
rect 31861 19873 31895 19907
rect 31895 19873 31904 19907
rect 31852 19864 31904 19873
rect 29092 19796 29144 19848
rect 29552 19796 29604 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 15844 19728 15896 19780
rect 18328 19728 18380 19780
rect 18880 19771 18932 19780
rect 18880 19737 18889 19771
rect 18889 19737 18923 19771
rect 18923 19737 18932 19771
rect 18880 19728 18932 19737
rect 19432 19728 19484 19780
rect 15936 19660 15988 19712
rect 16672 19660 16724 19712
rect 17132 19660 17184 19712
rect 17960 19660 18012 19712
rect 18788 19660 18840 19712
rect 22192 19728 22244 19780
rect 22652 19728 22704 19780
rect 19984 19660 20036 19712
rect 20720 19660 20772 19712
rect 23572 19660 23624 19712
rect 24124 19728 24176 19780
rect 30656 19728 30708 19780
rect 31576 19796 31628 19848
rect 37372 19796 37424 19848
rect 24492 19660 24544 19712
rect 29828 19703 29880 19712
rect 29828 19669 29837 19703
rect 29837 19669 29871 19703
rect 29871 19669 29880 19703
rect 29828 19660 29880 19669
rect 38108 19660 38160 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3056 19388 3108 19440
rect 3884 19388 3936 19440
rect 3976 19320 4028 19372
rect 11060 19388 11112 19440
rect 13452 19456 13504 19508
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 18328 19499 18380 19508
rect 18328 19465 18337 19499
rect 18337 19465 18371 19499
rect 18371 19465 18380 19499
rect 18328 19456 18380 19465
rect 21456 19456 21508 19508
rect 30104 19499 30156 19508
rect 15292 19388 15344 19440
rect 17224 19388 17276 19440
rect 17684 19431 17736 19440
rect 17684 19397 17693 19431
rect 17693 19397 17727 19431
rect 17727 19397 17736 19431
rect 17684 19388 17736 19397
rect 19340 19388 19392 19440
rect 20168 19388 20220 19440
rect 20812 19388 20864 19440
rect 3608 19252 3660 19304
rect 3792 19295 3844 19304
rect 3792 19261 3801 19295
rect 3801 19261 3835 19295
rect 3835 19261 3844 19295
rect 3792 19252 3844 19261
rect 10232 19363 10284 19372
rect 10232 19329 10241 19363
rect 10241 19329 10275 19363
rect 10275 19329 10284 19363
rect 10232 19320 10284 19329
rect 10324 19252 10376 19304
rect 10784 19252 10836 19304
rect 11152 19252 11204 19304
rect 16028 19320 16080 19372
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 20720 19363 20772 19372
rect 20720 19329 20729 19363
rect 20729 19329 20763 19363
rect 20763 19329 20772 19363
rect 20720 19320 20772 19329
rect 24032 19388 24084 19440
rect 30104 19465 30113 19499
rect 30113 19465 30147 19499
rect 30147 19465 30156 19499
rect 30104 19456 30156 19465
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 24492 19363 24544 19372
rect 24492 19329 24501 19363
rect 24501 19329 24535 19363
rect 24535 19329 24544 19363
rect 25780 19363 25832 19372
rect 24492 19320 24544 19329
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 25964 19363 26016 19372
rect 25964 19329 25973 19363
rect 25973 19329 26007 19363
rect 26007 19329 26016 19363
rect 25964 19320 26016 19329
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 20812 19295 20864 19304
rect 9864 19184 9916 19236
rect 15016 19184 15068 19236
rect 18052 19184 18104 19236
rect 10140 19116 10192 19168
rect 13452 19116 13504 19168
rect 13636 19116 13688 19168
rect 18696 19116 18748 19168
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 21180 19252 21232 19304
rect 23204 19295 23256 19304
rect 23204 19261 23213 19295
rect 23213 19261 23247 19295
rect 23247 19261 23256 19295
rect 23204 19252 23256 19261
rect 23664 19252 23716 19304
rect 23756 19184 23808 19236
rect 29828 19388 29880 19440
rect 27620 19320 27672 19372
rect 27988 19252 28040 19304
rect 30656 19320 30708 19372
rect 30932 19252 30984 19304
rect 26240 19184 26292 19236
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 30472 19116 30524 19168
rect 38292 19116 38344 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 9864 18912 9916 18964
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 10324 18955 10376 18964
rect 10324 18921 10333 18955
rect 10333 18921 10367 18955
rect 10367 18921 10376 18955
rect 10324 18912 10376 18921
rect 11980 18912 12032 18964
rect 13452 18912 13504 18964
rect 10692 18844 10744 18896
rect 2504 18776 2556 18828
rect 3332 18776 3384 18828
rect 4804 18819 4856 18828
rect 4804 18785 4813 18819
rect 4813 18785 4847 18819
rect 4847 18785 4856 18819
rect 4804 18776 4856 18785
rect 8852 18776 8904 18828
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 10140 18776 10192 18828
rect 10232 18708 10284 18760
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 11060 18751 11112 18760
rect 11060 18717 11094 18751
rect 11094 18717 11112 18751
rect 11060 18708 11112 18717
rect 2964 18640 3016 18692
rect 3332 18683 3384 18692
rect 3332 18649 3341 18683
rect 3341 18649 3375 18683
rect 3375 18649 3384 18683
rect 3332 18640 3384 18649
rect 3976 18683 4028 18692
rect 3976 18649 3985 18683
rect 3985 18649 4019 18683
rect 4019 18649 4028 18683
rect 3976 18640 4028 18649
rect 2228 18572 2280 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9588 18640 9640 18692
rect 13636 18844 13688 18896
rect 17224 18912 17276 18964
rect 20168 18955 20220 18964
rect 20168 18921 20177 18955
rect 20177 18921 20211 18955
rect 20211 18921 20220 18955
rect 20168 18912 20220 18921
rect 20812 18912 20864 18964
rect 31852 18912 31904 18964
rect 22376 18844 22428 18896
rect 22468 18844 22520 18896
rect 27436 18887 27488 18896
rect 27436 18853 27445 18887
rect 27445 18853 27479 18887
rect 27479 18853 27488 18887
rect 27436 18844 27488 18853
rect 28080 18844 28132 18896
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 22744 18776 22796 18828
rect 25964 18776 26016 18828
rect 28264 18819 28316 18828
rect 28264 18785 28273 18819
rect 28273 18785 28307 18819
rect 28307 18785 28316 18819
rect 28264 18776 28316 18785
rect 30656 18844 30708 18896
rect 37832 18819 37884 18828
rect 13544 18708 13596 18760
rect 13820 18708 13872 18760
rect 14556 18683 14608 18692
rect 14556 18649 14590 18683
rect 14590 18649 14608 18683
rect 14556 18640 14608 18649
rect 15200 18572 15252 18624
rect 16304 18708 16356 18760
rect 15752 18572 15804 18624
rect 17132 18572 17184 18624
rect 17316 18572 17368 18624
rect 17408 18572 17460 18624
rect 17592 18572 17644 18624
rect 20352 18708 20404 18760
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 21088 18708 21140 18760
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 23204 18708 23256 18760
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 27620 18751 27672 18760
rect 27620 18717 27629 18751
rect 27629 18717 27663 18751
rect 27663 18717 27672 18751
rect 27620 18708 27672 18717
rect 28448 18751 28500 18760
rect 28448 18717 28457 18751
rect 28457 18717 28491 18751
rect 28491 18717 28500 18751
rect 28448 18708 28500 18717
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 31668 18751 31720 18760
rect 28540 18708 28592 18717
rect 31668 18717 31677 18751
rect 31677 18717 31711 18751
rect 31711 18717 31720 18751
rect 31668 18708 31720 18717
rect 37832 18785 37841 18819
rect 37841 18785 37875 18819
rect 37875 18785 37884 18819
rect 37832 18776 37884 18785
rect 38108 18819 38160 18828
rect 38108 18785 38117 18819
rect 38117 18785 38151 18819
rect 38151 18785 38160 18819
rect 38108 18776 38160 18785
rect 38292 18819 38344 18828
rect 38292 18785 38301 18819
rect 38301 18785 38335 18819
rect 38335 18785 38344 18819
rect 38292 18776 38344 18785
rect 32496 18708 32548 18760
rect 17868 18640 17920 18692
rect 22376 18683 22428 18692
rect 20812 18615 20864 18624
rect 20812 18581 20821 18615
rect 20821 18581 20855 18615
rect 20855 18581 20864 18615
rect 20812 18572 20864 18581
rect 22376 18649 22385 18683
rect 22385 18649 22419 18683
rect 22419 18649 22428 18683
rect 22376 18640 22428 18649
rect 23848 18640 23900 18692
rect 30472 18640 30524 18692
rect 23204 18615 23256 18624
rect 23204 18581 23213 18615
rect 23213 18581 23247 18615
rect 23247 18581 23256 18615
rect 23204 18572 23256 18581
rect 24124 18572 24176 18624
rect 28264 18615 28316 18624
rect 28264 18581 28273 18615
rect 28273 18581 28307 18615
rect 28307 18581 28316 18615
rect 28264 18572 28316 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 11152 18368 11204 18420
rect 12348 18411 12400 18420
rect 12348 18377 12357 18411
rect 12357 18377 12391 18411
rect 12391 18377 12400 18411
rect 12348 18368 12400 18377
rect 16120 18368 16172 18420
rect 4620 18300 4672 18352
rect 3976 18232 4028 18284
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 9128 18232 9180 18284
rect 9588 18275 9640 18284
rect 9588 18241 9597 18275
rect 9597 18241 9631 18275
rect 9631 18241 9640 18275
rect 9588 18232 9640 18241
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 12164 18300 12216 18352
rect 16580 18300 16632 18352
rect 17684 18368 17736 18420
rect 20628 18411 20680 18420
rect 20628 18377 20637 18411
rect 20637 18377 20671 18411
rect 20671 18377 20680 18411
rect 20628 18368 20680 18377
rect 22468 18368 22520 18420
rect 22744 18368 22796 18420
rect 17224 18343 17276 18352
rect 17224 18309 17233 18343
rect 17233 18309 17267 18343
rect 17267 18309 17276 18343
rect 17224 18300 17276 18309
rect 11796 18232 11848 18284
rect 12440 18232 12492 18284
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 1860 18207 1912 18216
rect 1860 18173 1869 18207
rect 1869 18173 1903 18207
rect 1903 18173 1912 18207
rect 1860 18164 1912 18173
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 9680 18164 9732 18216
rect 15016 18164 15068 18216
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 16672 18232 16724 18284
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 18144 18300 18196 18352
rect 18420 18300 18472 18352
rect 20996 18300 21048 18352
rect 25780 18343 25832 18352
rect 16764 18164 16816 18216
rect 17592 18232 17644 18284
rect 20812 18232 20864 18284
rect 25780 18309 25789 18343
rect 25789 18309 25823 18343
rect 25823 18309 25832 18343
rect 25780 18300 25832 18309
rect 25872 18300 25924 18352
rect 26056 18300 26108 18352
rect 18236 18164 18288 18216
rect 21180 18164 21232 18216
rect 15844 18139 15896 18148
rect 15844 18105 15853 18139
rect 15853 18105 15887 18139
rect 15887 18105 15896 18139
rect 15844 18096 15896 18105
rect 17132 18096 17184 18148
rect 17316 18096 17368 18148
rect 9864 18028 9916 18080
rect 12992 18028 13044 18080
rect 13728 18028 13780 18080
rect 17592 18028 17644 18080
rect 18512 18096 18564 18148
rect 23480 18275 23532 18284
rect 23480 18241 23489 18275
rect 23489 18241 23523 18275
rect 23523 18241 23532 18275
rect 23664 18275 23716 18284
rect 23480 18232 23532 18241
rect 23664 18241 23673 18275
rect 23673 18241 23707 18275
rect 23707 18241 23716 18275
rect 23664 18232 23716 18241
rect 26516 18232 26568 18284
rect 28172 18368 28224 18420
rect 31668 18411 31720 18420
rect 31668 18377 31677 18411
rect 31677 18377 31711 18411
rect 31711 18377 31720 18411
rect 31668 18368 31720 18377
rect 30380 18300 30432 18352
rect 27436 18275 27488 18284
rect 27436 18241 27445 18275
rect 27445 18241 27479 18275
rect 27479 18241 27488 18275
rect 27436 18232 27488 18241
rect 27804 18232 27856 18284
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 27160 18164 27212 18216
rect 30472 18275 30524 18284
rect 21088 18028 21140 18080
rect 23572 18071 23624 18080
rect 23572 18037 23581 18071
rect 23581 18037 23615 18071
rect 23615 18037 23624 18071
rect 23572 18028 23624 18037
rect 25964 18028 26016 18080
rect 27160 18028 27212 18080
rect 30472 18241 30481 18275
rect 30481 18241 30515 18275
rect 30515 18241 30524 18275
rect 30472 18232 30524 18241
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 31484 18232 31536 18284
rect 32036 18232 32088 18284
rect 32496 18275 32548 18284
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 31116 18071 31168 18080
rect 31116 18037 31125 18071
rect 31125 18037 31159 18071
rect 31159 18037 31168 18071
rect 31116 18028 31168 18037
rect 31208 18028 31260 18080
rect 36452 18028 36504 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1860 17824 1912 17876
rect 2044 17824 2096 17876
rect 9128 17824 9180 17876
rect 13084 17867 13136 17876
rect 13084 17833 13093 17867
rect 13093 17833 13127 17867
rect 13127 17833 13136 17867
rect 13084 17824 13136 17833
rect 14556 17867 14608 17876
rect 14556 17833 14565 17867
rect 14565 17833 14599 17867
rect 14599 17833 14608 17867
rect 14556 17824 14608 17833
rect 18144 17867 18196 17876
rect 18144 17833 18153 17867
rect 18153 17833 18187 17867
rect 18187 17833 18196 17867
rect 18144 17824 18196 17833
rect 3608 17688 3660 17740
rect 4804 17688 4856 17740
rect 9680 17688 9732 17740
rect 3240 17620 3292 17672
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 4712 17620 4764 17672
rect 8852 17620 8904 17672
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 10416 17620 10468 17672
rect 10784 17620 10836 17672
rect 13820 17620 13872 17672
rect 15568 17756 15620 17808
rect 16212 17756 16264 17808
rect 23112 17824 23164 17876
rect 27436 17824 27488 17876
rect 27804 17824 27856 17876
rect 30472 17824 30524 17876
rect 32036 17867 32088 17876
rect 20352 17799 20404 17808
rect 20352 17765 20361 17799
rect 20361 17765 20395 17799
rect 20395 17765 20404 17799
rect 20352 17756 20404 17765
rect 16672 17688 16724 17740
rect 17316 17688 17368 17740
rect 19156 17688 19208 17740
rect 21180 17688 21232 17740
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15200 17663 15252 17672
rect 15016 17620 15068 17629
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 20996 17620 21048 17672
rect 25964 17663 26016 17672
rect 16580 17552 16632 17604
rect 22100 17552 22152 17604
rect 23020 17552 23072 17604
rect 24952 17552 25004 17604
rect 25964 17629 25973 17663
rect 25973 17629 26007 17663
rect 26007 17629 26016 17663
rect 25964 17620 26016 17629
rect 26332 17663 26384 17672
rect 26332 17629 26341 17663
rect 26341 17629 26375 17663
rect 26375 17629 26384 17663
rect 26332 17620 26384 17629
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 27160 17620 27212 17672
rect 28632 17756 28684 17808
rect 29000 17756 29052 17808
rect 31208 17756 31260 17808
rect 32036 17833 32045 17867
rect 32045 17833 32079 17867
rect 32079 17833 32088 17867
rect 32036 17824 32088 17833
rect 28264 17663 28316 17672
rect 28264 17629 28273 17663
rect 28273 17629 28307 17663
rect 28307 17629 28316 17663
rect 28264 17620 28316 17629
rect 28448 17620 28500 17672
rect 31116 17688 31168 17740
rect 36452 17731 36504 17740
rect 36452 17697 36461 17731
rect 36461 17697 36495 17731
rect 36495 17697 36504 17731
rect 36452 17688 36504 17697
rect 38292 17731 38344 17740
rect 38292 17697 38301 17731
rect 38301 17697 38335 17731
rect 38335 17697 38344 17731
rect 38292 17688 38344 17697
rect 30748 17663 30800 17672
rect 30748 17629 30757 17663
rect 30757 17629 30791 17663
rect 30791 17629 30800 17663
rect 30748 17620 30800 17629
rect 25688 17552 25740 17604
rect 3516 17484 3568 17536
rect 14924 17484 14976 17536
rect 16856 17484 16908 17536
rect 17592 17484 17644 17536
rect 22008 17484 22060 17536
rect 23112 17484 23164 17536
rect 26148 17595 26200 17604
rect 26148 17561 26157 17595
rect 26157 17561 26191 17595
rect 26191 17561 26200 17595
rect 31484 17620 31536 17672
rect 26148 17552 26200 17561
rect 31024 17552 31076 17604
rect 37556 17552 37608 17604
rect 27160 17484 27212 17536
rect 28540 17484 28592 17536
rect 30288 17484 30340 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 3240 17280 3292 17332
rect 3516 17255 3568 17264
rect 3516 17221 3525 17255
rect 3525 17221 3559 17255
rect 3559 17221 3568 17255
rect 3516 17212 3568 17221
rect 12624 17212 12676 17264
rect 13544 17212 13596 17264
rect 16948 17212 17000 17264
rect 17316 17255 17368 17264
rect 17316 17221 17325 17255
rect 17325 17221 17359 17255
rect 17359 17221 17368 17255
rect 17316 17212 17368 17221
rect 17776 17212 17828 17264
rect 21088 17255 21140 17264
rect 21088 17221 21097 17255
rect 21097 17221 21131 17255
rect 21131 17221 21140 17255
rect 21088 17212 21140 17221
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13636 17144 13688 17196
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 14648 17144 14700 17196
rect 16028 17187 16080 17196
rect 16028 17153 16062 17187
rect 16062 17153 16080 17187
rect 17500 17187 17552 17196
rect 16028 17144 16080 17153
rect 1860 17119 1912 17128
rect 1860 17085 1869 17119
rect 1869 17085 1903 17119
rect 1903 17085 1912 17119
rect 1860 17076 1912 17085
rect 2136 17076 2188 17128
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 20996 17187 21048 17196
rect 19340 17076 19392 17128
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 12900 17008 12952 17060
rect 13176 17051 13228 17060
rect 13176 17017 13185 17051
rect 13185 17017 13219 17051
rect 13219 17017 13228 17051
rect 13176 17008 13228 17017
rect 14188 16940 14240 16992
rect 14464 16940 14516 16992
rect 17040 17008 17092 17060
rect 19984 17008 20036 17060
rect 23204 17280 23256 17332
rect 23664 17280 23716 17332
rect 26056 17280 26108 17332
rect 23112 17255 23164 17264
rect 23112 17221 23121 17255
rect 23121 17221 23155 17255
rect 23155 17221 23164 17255
rect 23112 17212 23164 17221
rect 22376 17144 22428 17196
rect 23020 17144 23072 17196
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 26332 17280 26384 17332
rect 30288 17323 30340 17332
rect 30288 17289 30297 17323
rect 30297 17289 30331 17323
rect 30331 17289 30340 17323
rect 30288 17280 30340 17289
rect 37556 17323 37608 17332
rect 37556 17289 37565 17323
rect 37565 17289 37599 17323
rect 37599 17289 37608 17323
rect 37556 17280 37608 17289
rect 23296 17144 23348 17153
rect 23388 17076 23440 17128
rect 23572 17008 23624 17060
rect 15292 16940 15344 16992
rect 16212 16983 16264 16992
rect 16212 16949 16221 16983
rect 16221 16949 16255 16983
rect 16255 16949 16264 16983
rect 16212 16940 16264 16949
rect 16948 16940 17000 16992
rect 17960 16940 18012 16992
rect 23020 16940 23072 16992
rect 23756 16940 23808 16992
rect 25320 17119 25372 17128
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 26056 17076 26108 17128
rect 27160 17187 27212 17196
rect 27160 17153 27169 17187
rect 27169 17153 27203 17187
rect 27203 17153 27212 17187
rect 27160 17144 27212 17153
rect 27436 17187 27488 17196
rect 27436 17153 27445 17187
rect 27445 17153 27479 17187
rect 27479 17153 27488 17187
rect 27436 17144 27488 17153
rect 30104 17187 30156 17196
rect 30104 17153 30113 17187
rect 30113 17153 30147 17187
rect 30147 17153 30156 17187
rect 30104 17144 30156 17153
rect 30380 17187 30432 17196
rect 30380 17153 30389 17187
rect 30389 17153 30423 17187
rect 30423 17153 30432 17187
rect 30380 17144 30432 17153
rect 37280 17144 37332 17196
rect 38016 17144 38068 17196
rect 26240 17076 26292 17128
rect 27620 17076 27672 17128
rect 33876 17008 33928 17060
rect 25964 16983 26016 16992
rect 25964 16949 25973 16983
rect 25973 16949 26007 16983
rect 26007 16949 26016 16983
rect 25964 16940 26016 16949
rect 26148 16940 26200 16992
rect 27344 16983 27396 16992
rect 27344 16949 27353 16983
rect 27353 16949 27387 16983
rect 27387 16949 27396 16983
rect 27344 16940 27396 16949
rect 28356 16940 28408 16992
rect 36636 16940 36688 16992
rect 38108 16983 38160 16992
rect 38108 16949 38117 16983
rect 38117 16949 38151 16983
rect 38151 16949 38160 16983
rect 38108 16940 38160 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2136 16779 2188 16788
rect 2136 16745 2145 16779
rect 2145 16745 2179 16779
rect 2179 16745 2188 16779
rect 2136 16736 2188 16745
rect 3792 16736 3844 16788
rect 3976 16736 4028 16788
rect 12900 16779 12952 16788
rect 9128 16600 9180 16652
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 8852 16532 8904 16584
rect 10232 16532 10284 16584
rect 12624 16668 12676 16720
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 13176 16736 13228 16788
rect 13636 16736 13688 16788
rect 14464 16736 14516 16788
rect 14648 16736 14700 16788
rect 16764 16736 16816 16788
rect 17408 16736 17460 16788
rect 17684 16779 17736 16788
rect 17684 16745 17693 16779
rect 17693 16745 17727 16779
rect 17727 16745 17736 16779
rect 17684 16736 17736 16745
rect 27620 16736 27672 16788
rect 30380 16736 30432 16788
rect 2964 16396 3016 16448
rect 4804 16464 4856 16516
rect 12440 16532 12492 16584
rect 13360 16575 13412 16584
rect 8484 16396 8536 16448
rect 11796 16464 11848 16516
rect 12624 16507 12676 16516
rect 12624 16473 12633 16507
rect 12633 16473 12667 16507
rect 12667 16473 12676 16507
rect 12624 16464 12676 16473
rect 11428 16439 11480 16448
rect 11428 16405 11437 16439
rect 11437 16405 11471 16439
rect 11471 16405 11480 16439
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 14188 16600 14240 16652
rect 15292 16532 15344 16584
rect 16856 16600 16908 16652
rect 25872 16600 25924 16652
rect 25964 16600 26016 16652
rect 27620 16600 27672 16652
rect 28356 16643 28408 16652
rect 28356 16609 28365 16643
rect 28365 16609 28399 16643
rect 28399 16609 28408 16643
rect 28356 16600 28408 16609
rect 30472 16668 30524 16720
rect 38016 16736 38068 16788
rect 38108 16668 38160 16720
rect 36636 16643 36688 16652
rect 36636 16609 36645 16643
rect 36645 16609 36679 16643
rect 36679 16609 36688 16643
rect 36636 16600 36688 16609
rect 38292 16643 38344 16652
rect 38292 16609 38301 16643
rect 38301 16609 38335 16643
rect 38335 16609 38344 16643
rect 38292 16600 38344 16609
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 17592 16575 17644 16584
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 17684 16532 17736 16584
rect 18512 16532 18564 16584
rect 21732 16532 21784 16584
rect 23296 16532 23348 16584
rect 28264 16575 28316 16584
rect 28264 16541 28273 16575
rect 28273 16541 28307 16575
rect 28307 16541 28316 16575
rect 28264 16532 28316 16541
rect 30932 16532 30984 16584
rect 31300 16575 31352 16584
rect 31300 16541 31309 16575
rect 31309 16541 31343 16575
rect 31343 16541 31352 16575
rect 31300 16532 31352 16541
rect 15660 16439 15712 16448
rect 11428 16396 11480 16405
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 21272 16396 21324 16448
rect 21824 16396 21876 16448
rect 23756 16396 23808 16448
rect 24308 16396 24360 16448
rect 27896 16439 27948 16448
rect 27896 16405 27905 16439
rect 27905 16405 27939 16439
rect 27939 16405 27948 16439
rect 27896 16396 27948 16405
rect 30104 16396 30156 16448
rect 30288 16396 30340 16448
rect 37372 16396 37424 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 12440 16192 12492 16244
rect 12808 16192 12860 16244
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 3240 16124 3292 16176
rect 3700 16124 3752 16176
rect 17224 16192 17276 16244
rect 23296 16192 23348 16244
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 4436 16056 4488 16108
rect 4620 16056 4672 16108
rect 10232 16056 10284 16108
rect 10508 16031 10560 16040
rect 5632 15920 5684 15972
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 10508 15988 10560 15997
rect 11796 15988 11848 16040
rect 11520 15920 11572 15972
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 17316 16056 17368 16108
rect 18604 16124 18656 16176
rect 17960 16056 18012 16108
rect 14924 15988 14976 16040
rect 10508 15852 10560 15904
rect 12716 15852 12768 15904
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 30288 16124 30340 16176
rect 21272 16099 21324 16108
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 25320 16056 25372 16108
rect 27620 16099 27672 16108
rect 27620 16065 27629 16099
rect 27629 16065 27663 16099
rect 27663 16065 27672 16099
rect 27620 16056 27672 16065
rect 23572 15988 23624 16040
rect 27436 15988 27488 16040
rect 27252 15920 27304 15972
rect 30104 16056 30156 16108
rect 31300 16099 31352 16108
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 37740 16056 37792 16108
rect 28264 15920 28316 15972
rect 30012 15988 30064 16040
rect 30380 15988 30432 16040
rect 30932 15920 30984 15972
rect 19248 15895 19300 15904
rect 19248 15861 19257 15895
rect 19257 15861 19291 15895
rect 19291 15861 19300 15895
rect 19248 15852 19300 15861
rect 28724 15895 28776 15904
rect 28724 15861 28733 15895
rect 28733 15861 28767 15895
rect 28767 15861 28776 15895
rect 28724 15852 28776 15861
rect 30196 15852 30248 15904
rect 36636 15852 36688 15904
rect 37648 15895 37700 15904
rect 37648 15861 37657 15895
rect 37657 15861 37691 15895
rect 37691 15861 37700 15895
rect 37648 15852 37700 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4528 15648 4580 15700
rect 4712 15648 4764 15700
rect 11428 15648 11480 15700
rect 11520 15648 11572 15700
rect 37464 15648 37516 15700
rect 2228 15580 2280 15632
rect 2872 15555 2924 15564
rect 2872 15521 2881 15555
rect 2881 15521 2915 15555
rect 2915 15521 2924 15555
rect 2872 15512 2924 15521
rect 10324 15512 10376 15564
rect 17960 15623 18012 15632
rect 17960 15589 17969 15623
rect 17969 15589 18003 15623
rect 18003 15589 18012 15623
rect 17960 15580 18012 15589
rect 23204 15623 23256 15632
rect 23204 15589 23213 15623
rect 23213 15589 23247 15623
rect 23247 15589 23256 15623
rect 23204 15580 23256 15589
rect 27988 15580 28040 15632
rect 30564 15623 30616 15632
rect 14924 15555 14976 15564
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 9588 15487 9640 15496
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 3240 15419 3292 15428
rect 3240 15385 3249 15419
rect 3249 15385 3283 15419
rect 3283 15385 3292 15419
rect 3240 15376 3292 15385
rect 2320 15308 2372 15360
rect 4712 15376 4764 15428
rect 13728 15444 13780 15496
rect 15476 15444 15528 15496
rect 16212 15444 16264 15496
rect 18236 15512 18288 15564
rect 18696 15512 18748 15564
rect 13544 15376 13596 15428
rect 17040 15376 17092 15428
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 19248 15444 19300 15496
rect 23572 15512 23624 15564
rect 26700 15555 26752 15564
rect 26700 15521 26709 15555
rect 26709 15521 26743 15555
rect 26743 15521 26752 15555
rect 27436 15555 27488 15564
rect 26700 15512 26752 15521
rect 27436 15521 27445 15555
rect 27445 15521 27479 15555
rect 27479 15521 27488 15555
rect 27436 15512 27488 15521
rect 27252 15444 27304 15496
rect 29092 15512 29144 15564
rect 30564 15589 30573 15623
rect 30573 15589 30607 15623
rect 30607 15589 30616 15623
rect 30564 15580 30616 15589
rect 37648 15580 37700 15632
rect 36636 15555 36688 15564
rect 36636 15521 36645 15555
rect 36645 15521 36679 15555
rect 36679 15521 36688 15555
rect 36636 15512 36688 15521
rect 38292 15555 38344 15564
rect 38292 15521 38301 15555
rect 38301 15521 38335 15555
rect 38335 15521 38344 15555
rect 38292 15512 38344 15521
rect 30380 15444 30432 15496
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 30656 15444 30708 15453
rect 20076 15376 20128 15428
rect 4804 15308 4856 15360
rect 9772 15308 9824 15360
rect 12440 15308 12492 15360
rect 16488 15308 16540 15360
rect 17592 15308 17644 15360
rect 20168 15308 20220 15360
rect 25872 15308 25924 15360
rect 28264 15308 28316 15360
rect 30104 15308 30156 15360
rect 30840 15308 30892 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 13360 15104 13412 15156
rect 19156 15104 19208 15156
rect 19984 15104 20036 15156
rect 20076 15147 20128 15156
rect 20076 15113 20085 15147
rect 20085 15113 20119 15147
rect 20119 15113 20128 15147
rect 20076 15104 20128 15113
rect 21916 15104 21968 15156
rect 23572 15147 23624 15156
rect 23572 15113 23581 15147
rect 23581 15113 23615 15147
rect 23615 15113 23624 15147
rect 23572 15104 23624 15113
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 13268 14968 13320 15020
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 14188 14968 14240 15020
rect 21272 15036 21324 15088
rect 30656 15147 30708 15156
rect 30656 15113 30665 15147
rect 30665 15113 30699 15147
rect 30699 15113 30708 15147
rect 30656 15104 30708 15113
rect 26700 15036 26752 15088
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 12532 14943 12584 14952
rect 2780 14900 2832 14909
rect 12532 14909 12549 14943
rect 12549 14909 12583 14943
rect 12583 14909 12584 14943
rect 12532 14900 12584 14909
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 14648 14832 14700 14884
rect 16120 14832 16172 14884
rect 19984 15011 20036 15020
rect 19984 14977 20026 15011
rect 20026 14977 20036 15011
rect 21088 15011 21140 15020
rect 19984 14968 20036 14977
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 24952 15011 25004 15020
rect 24952 14977 24961 15011
rect 24961 14977 24995 15011
rect 24995 14977 25004 15011
rect 24952 14968 25004 14977
rect 27252 14968 27304 15020
rect 30288 15011 30340 15020
rect 30288 14977 30297 15011
rect 30297 14977 30331 15011
rect 30331 14977 30340 15011
rect 30288 14968 30340 14977
rect 12808 14764 12860 14816
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 22836 14832 22888 14884
rect 20996 14764 21048 14816
rect 21272 14764 21324 14816
rect 29092 14900 29144 14952
rect 30196 14943 30248 14952
rect 30196 14909 30205 14943
rect 30205 14909 30239 14943
rect 30239 14909 30248 14943
rect 30196 14900 30248 14909
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 3240 14560 3292 14612
rect 16672 14560 16724 14612
rect 18420 14560 18472 14612
rect 19984 14560 20036 14612
rect 21088 14560 21140 14612
rect 27252 14603 27304 14612
rect 27252 14569 27261 14603
rect 27261 14569 27295 14603
rect 27295 14569 27304 14603
rect 27252 14560 27304 14569
rect 27620 14560 27672 14612
rect 29000 14560 29052 14612
rect 22376 14535 22428 14544
rect 22376 14501 22385 14535
rect 22385 14501 22419 14535
rect 22419 14501 22428 14535
rect 22376 14492 22428 14501
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 3056 14356 3108 14408
rect 10416 14356 10468 14408
rect 14924 14356 14976 14408
rect 22008 14424 22060 14476
rect 16304 14356 16356 14408
rect 10232 14288 10284 14340
rect 14096 14288 14148 14340
rect 16212 14288 16264 14340
rect 19432 14356 19484 14408
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 27436 14399 27488 14408
rect 22100 14356 22152 14365
rect 27436 14365 27442 14399
rect 27442 14365 27476 14399
rect 27476 14365 27488 14399
rect 27436 14356 27488 14365
rect 27896 14399 27948 14408
rect 27896 14365 27905 14399
rect 27905 14365 27939 14399
rect 27939 14365 27948 14399
rect 27896 14356 27948 14365
rect 21824 14288 21876 14340
rect 24860 14288 24912 14340
rect 26516 14288 26568 14340
rect 29828 14288 29880 14340
rect 2872 14220 2924 14272
rect 12716 14220 12768 14272
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 17592 14220 17644 14272
rect 20076 14220 20128 14272
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 26332 14220 26384 14272
rect 30104 14220 30156 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2228 14059 2280 14068
rect 2228 14025 2237 14059
rect 2237 14025 2271 14059
rect 2271 14025 2280 14059
rect 2228 14016 2280 14025
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 12624 14059 12676 14068
rect 12624 14025 12633 14059
rect 12633 14025 12667 14059
rect 12667 14025 12676 14059
rect 12624 14016 12676 14025
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 16304 14016 16356 14068
rect 19432 14016 19484 14068
rect 19984 14016 20036 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 3148 13880 3200 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 13544 13880 13596 13932
rect 14648 13880 14700 13932
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 15568 13880 15620 13932
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 16948 13880 17000 13932
rect 17224 13880 17276 13932
rect 19248 13948 19300 14000
rect 25688 14016 25740 14068
rect 27896 14059 27948 14068
rect 27896 14025 27905 14059
rect 27905 14025 27939 14059
rect 27939 14025 27948 14059
rect 27896 14016 27948 14025
rect 22008 13948 22060 14000
rect 19156 13880 19208 13932
rect 14740 13812 14792 13821
rect 16488 13812 16540 13864
rect 22376 13880 22428 13932
rect 24952 13948 25004 14000
rect 25136 13880 25188 13932
rect 27988 13880 28040 13932
rect 29184 13923 29236 13932
rect 29184 13889 29193 13923
rect 29193 13889 29227 13923
rect 29227 13889 29236 13923
rect 29184 13880 29236 13889
rect 29828 13923 29880 13932
rect 29828 13889 29837 13923
rect 29837 13889 29871 13923
rect 29871 13889 29880 13923
rect 29828 13880 29880 13889
rect 30104 13923 30156 13932
rect 30104 13889 30113 13923
rect 30113 13889 30147 13923
rect 30147 13889 30156 13923
rect 30104 13880 30156 13889
rect 9128 13744 9180 13796
rect 12624 13744 12676 13796
rect 16672 13744 16724 13796
rect 18420 13676 18472 13728
rect 28080 13812 28132 13864
rect 28724 13812 28776 13864
rect 29920 13812 29972 13864
rect 22744 13676 22796 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10048 13472 10100 13524
rect 10324 13472 10376 13524
rect 13268 13472 13320 13524
rect 14740 13472 14792 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 18512 13472 18564 13524
rect 21916 13515 21968 13524
rect 21916 13481 21925 13515
rect 21925 13481 21959 13515
rect 21959 13481 21968 13515
rect 21916 13472 21968 13481
rect 12532 13404 12584 13456
rect 12808 13404 12860 13456
rect 16672 13404 16724 13456
rect 10416 13379 10468 13388
rect 10416 13345 10425 13379
rect 10425 13345 10459 13379
rect 10459 13345 10468 13379
rect 10416 13336 10468 13345
rect 17960 13336 18012 13388
rect 22192 13472 22244 13524
rect 23756 13515 23808 13524
rect 23756 13481 23765 13515
rect 23765 13481 23799 13515
rect 23799 13481 23808 13515
rect 23756 13472 23808 13481
rect 25136 13515 25188 13524
rect 25136 13481 25145 13515
rect 25145 13481 25179 13515
rect 25179 13481 25188 13515
rect 25136 13472 25188 13481
rect 25688 13472 25740 13524
rect 11244 13268 11296 13320
rect 12256 13268 12308 13320
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17500 13268 17552 13320
rect 21824 13268 21876 13320
rect 22744 13311 22796 13320
rect 9496 13200 9548 13252
rect 10416 13200 10468 13252
rect 10692 13243 10744 13252
rect 10692 13209 10726 13243
rect 10726 13209 10744 13243
rect 10692 13200 10744 13209
rect 14188 13200 14240 13252
rect 17776 13243 17828 13252
rect 17776 13209 17785 13243
rect 17785 13209 17819 13243
rect 17819 13209 17828 13243
rect 22744 13277 22753 13311
rect 22753 13277 22787 13311
rect 22787 13277 22796 13311
rect 22744 13268 22796 13277
rect 24860 13268 24912 13320
rect 27528 13472 27580 13524
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 27804 13311 27856 13320
rect 26792 13268 26844 13277
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 28080 13311 28132 13320
rect 28080 13277 28089 13311
rect 28089 13277 28123 13311
rect 28123 13277 28132 13311
rect 28080 13268 28132 13277
rect 38292 13268 38344 13320
rect 17776 13200 17828 13209
rect 29920 13200 29972 13252
rect 26332 13175 26384 13184
rect 26332 13141 26341 13175
rect 26341 13141 26375 13175
rect 26375 13141 26384 13175
rect 26332 13132 26384 13141
rect 27620 13175 27672 13184
rect 27620 13141 27629 13175
rect 27629 13141 27663 13175
rect 27663 13141 27672 13175
rect 27620 13132 27672 13141
rect 27988 13175 28040 13184
rect 27988 13141 27997 13175
rect 27997 13141 28031 13175
rect 28031 13141 28040 13175
rect 27988 13132 28040 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 14188 12928 14240 12980
rect 17500 12928 17552 12980
rect 17960 12971 18012 12980
rect 17960 12937 17969 12971
rect 17969 12937 18003 12971
rect 18003 12937 18012 12971
rect 17960 12928 18012 12937
rect 19248 12928 19300 12980
rect 20168 12928 20220 12980
rect 26792 12928 26844 12980
rect 27804 12971 27856 12980
rect 27804 12937 27813 12971
rect 27813 12937 27847 12971
rect 27847 12937 27856 12971
rect 27804 12928 27856 12937
rect 10692 12903 10744 12912
rect 10692 12869 10701 12903
rect 10701 12869 10735 12903
rect 10735 12869 10744 12903
rect 10692 12860 10744 12869
rect 14280 12860 14332 12912
rect 14648 12860 14700 12912
rect 2320 12792 2372 12844
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 10416 12792 10468 12844
rect 11244 12724 11296 12776
rect 12716 12724 12768 12776
rect 14004 12792 14056 12844
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 15660 12792 15712 12844
rect 16488 12860 16540 12912
rect 17592 12860 17644 12912
rect 17776 12860 17828 12912
rect 17408 12835 17460 12844
rect 4068 12656 4120 12708
rect 9956 12656 10008 12708
rect 16120 12724 16172 12776
rect 17408 12801 17417 12835
rect 17417 12801 17451 12835
rect 17451 12801 17460 12835
rect 17408 12792 17460 12801
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 18236 12835 18288 12844
rect 18236 12801 18245 12835
rect 18245 12801 18279 12835
rect 18279 12801 18288 12835
rect 18420 12835 18472 12844
rect 18236 12792 18288 12801
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 19248 12835 19300 12844
rect 13452 12656 13504 12708
rect 14556 12699 14608 12708
rect 14556 12665 14565 12699
rect 14565 12665 14599 12699
rect 14599 12665 14608 12699
rect 14556 12656 14608 12665
rect 15292 12656 15344 12708
rect 16212 12656 16264 12708
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 19432 12792 19484 12844
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 19340 12724 19392 12776
rect 29184 12860 29236 12912
rect 25688 12792 25740 12844
rect 27620 12792 27672 12844
rect 37924 12792 37976 12844
rect 27160 12724 27212 12776
rect 27436 12724 27488 12776
rect 1768 12588 1820 12640
rect 10508 12631 10560 12640
rect 10508 12597 10517 12631
rect 10517 12597 10551 12631
rect 10551 12597 10560 12631
rect 10508 12588 10560 12597
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 13268 12588 13320 12640
rect 15752 12588 15804 12640
rect 17132 12588 17184 12640
rect 19156 12588 19208 12640
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 28080 12588 28132 12640
rect 38108 12588 38160 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10508 12384 10560 12436
rect 13360 12384 13412 12436
rect 13452 12384 13504 12436
rect 17316 12384 17368 12436
rect 18420 12384 18472 12436
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20536 12384 20588 12436
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22100 12384 22152 12393
rect 27988 12384 28040 12436
rect 14188 12316 14240 12368
rect 15568 12316 15620 12368
rect 17408 12316 17460 12368
rect 18144 12316 18196 12368
rect 1768 12291 1820 12300
rect 1768 12257 1777 12291
rect 1777 12257 1811 12291
rect 1811 12257 1820 12291
rect 1768 12248 1820 12257
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 10232 12248 10284 12300
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 10324 12180 10376 12232
rect 12348 12248 12400 12300
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 12900 12248 12952 12300
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12716 12180 12768 12232
rect 15660 12248 15712 12300
rect 15752 12248 15804 12300
rect 37188 12291 37240 12300
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 16120 12223 16172 12232
rect 14740 12180 14792 12189
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 17592 12180 17644 12232
rect 12532 12112 12584 12164
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12624 12044 12676 12096
rect 16212 12044 16264 12096
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 18420 12180 18472 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 37188 12257 37197 12291
rect 37197 12257 37231 12291
rect 37231 12257 37240 12291
rect 37188 12248 37240 12257
rect 38108 12291 38160 12300
rect 38108 12257 38117 12291
rect 38117 12257 38151 12291
rect 38151 12257 38160 12291
rect 38108 12248 38160 12257
rect 38292 12291 38344 12300
rect 38292 12257 38301 12291
rect 38301 12257 38335 12291
rect 38335 12257 38344 12291
rect 38292 12248 38344 12257
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20904 12223 20956 12232
rect 20260 12180 20312 12189
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 21456 12180 21508 12232
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 27804 12180 27856 12232
rect 28080 12223 28132 12232
rect 28080 12189 28089 12223
rect 28089 12189 28123 12223
rect 28123 12189 28132 12223
rect 28080 12180 28132 12189
rect 19432 12112 19484 12164
rect 20076 12112 20128 12164
rect 19340 12044 19392 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 12900 11840 12952 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 16120 11840 16172 11892
rect 17316 11840 17368 11892
rect 12532 11772 12584 11824
rect 1584 11704 1636 11756
rect 9772 11704 9824 11756
rect 10508 11704 10560 11756
rect 11980 11704 12032 11756
rect 11796 11611 11848 11620
rect 11796 11577 11805 11611
rect 11805 11577 11839 11611
rect 11839 11577 11848 11611
rect 11796 11568 11848 11577
rect 11612 11500 11664 11552
rect 12716 11500 12768 11552
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14648 11704 14700 11756
rect 14464 11568 14516 11620
rect 15752 11772 15804 11824
rect 18880 11772 18932 11824
rect 15568 11704 15620 11756
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 16212 11704 16264 11756
rect 17224 11636 17276 11688
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 18420 11679 18472 11688
rect 16396 11568 16448 11620
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 19340 11704 19392 11756
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 20076 11747 20128 11756
rect 19800 11704 19852 11713
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 20904 11704 20956 11756
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 21916 11840 21968 11892
rect 21548 11772 21600 11824
rect 22744 11772 22796 11824
rect 19156 11568 19208 11620
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 37372 11704 37424 11756
rect 20260 11636 20312 11645
rect 21456 11611 21508 11620
rect 21456 11577 21465 11611
rect 21465 11577 21499 11611
rect 21499 11577 21508 11611
rect 21456 11568 21508 11577
rect 16212 11500 16264 11552
rect 16304 11500 16356 11552
rect 20168 11500 20220 11552
rect 21180 11500 21232 11552
rect 21548 11500 21600 11552
rect 38108 11500 38160 11552
rect 38292 11543 38344 11552
rect 38292 11509 38301 11543
rect 38301 11509 38335 11543
rect 38335 11509 38344 11543
rect 38292 11500 38344 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12256 11339 12308 11348
rect 12256 11305 12265 11339
rect 12265 11305 12299 11339
rect 12299 11305 12308 11339
rect 12256 11296 12308 11305
rect 12348 11296 12400 11348
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 12900 11296 12952 11348
rect 15844 11296 15896 11348
rect 10508 11228 10560 11280
rect 18420 11296 18472 11348
rect 21180 11296 21232 11348
rect 17224 11228 17276 11280
rect 18512 11228 18564 11280
rect 21824 11228 21876 11280
rect 3056 11160 3108 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3240 11067 3292 11076
rect 3240 11033 3249 11067
rect 3249 11033 3283 11067
rect 3283 11033 3292 11067
rect 3240 11024 3292 11033
rect 16396 11160 16448 11212
rect 19800 11160 19852 11212
rect 37188 11203 37240 11212
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 20168 11092 20220 11144
rect 37188 11169 37197 11203
rect 37197 11169 37231 11203
rect 37231 11169 37240 11203
rect 37188 11160 37240 11169
rect 38108 11203 38160 11212
rect 38108 11169 38117 11203
rect 38117 11169 38151 11203
rect 38151 11169 38160 11203
rect 38108 11160 38160 11169
rect 38292 11203 38344 11212
rect 38292 11169 38301 11203
rect 38301 11169 38335 11203
rect 38335 11169 38344 11203
rect 38292 11160 38344 11169
rect 18328 11024 18380 11076
rect 16212 10956 16264 11008
rect 20812 10956 20864 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3240 10752 3292 10804
rect 2964 10616 3016 10668
rect 18328 10616 18380 10668
rect 3424 10548 3476 10600
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 18604 10208 18656 10260
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 32956 10004 33008 10056
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2872 9528 2924 9580
rect 23848 9571 23900 9580
rect 4712 9460 4764 9512
rect 23848 9537 23857 9571
rect 23857 9537 23891 9571
rect 23891 9537 23900 9571
rect 23848 9528 23900 9537
rect 34520 9460 34572 9512
rect 29092 9392 29144 9444
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 3240 9324 3292 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2044 9052 2096 9104
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 4712 8916 4764 8968
rect 34796 8916 34848 8968
rect 38292 8916 38344 8968
rect 1584 8891 1636 8900
rect 1584 8857 1593 8891
rect 1593 8857 1627 8891
rect 1627 8857 1636 8891
rect 1584 8848 1636 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 20352 8440 20404 8492
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 37832 8279 37884 8288
rect 37832 8245 37841 8279
rect 37841 8245 37875 8279
rect 37875 8245 37884 8279
rect 37832 8236 37884 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 37188 7939 37240 7948
rect 37188 7905 37197 7939
rect 37197 7905 37231 7939
rect 37231 7905 37240 7939
rect 37188 7896 37240 7905
rect 37832 7896 37884 7948
rect 37556 7760 37608 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 37556 7531 37608 7540
rect 37556 7497 37565 7531
rect 37565 7497 37599 7531
rect 37599 7497 37608 7531
rect 37556 7488 37608 7497
rect 37372 7352 37424 7404
rect 38016 7352 38068 7404
rect 3424 7148 3476 7200
rect 5356 7191 5408 7200
rect 5356 7157 5365 7191
rect 5365 7157 5399 7191
rect 5399 7157 5408 7191
rect 5356 7148 5408 7157
rect 38108 7148 38160 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 37188 6851 37240 6860
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 38108 6851 38160 6860
rect 38108 6817 38117 6851
rect 38117 6817 38151 6851
rect 38151 6817 38160 6851
rect 38108 6808 38160 6817
rect 38292 6851 38344 6860
rect 38292 6817 38301 6851
rect 38301 6817 38335 6851
rect 38335 6817 38344 6851
rect 38292 6808 38344 6817
rect 2412 6672 2464 6724
rect 5540 6715 5592 6724
rect 5540 6681 5549 6715
rect 5549 6681 5583 6715
rect 5583 6681 5592 6715
rect 5540 6672 5592 6681
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 4712 6332 4764 6384
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 4068 6264 4120 6316
rect 37280 6264 37332 6316
rect 38108 6060 38160 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 39304 5788 39356 5840
rect 38108 5763 38160 5772
rect 38108 5729 38117 5763
rect 38117 5729 38151 5763
rect 38151 5729 38160 5763
rect 38108 5720 38160 5729
rect 1860 5652 1912 5704
rect 3148 5652 3200 5704
rect 3608 5652 3660 5704
rect 20812 5652 20864 5704
rect 38292 5695 38344 5704
rect 38292 5661 38301 5695
rect 38301 5661 38335 5695
rect 38335 5661 38344 5695
rect 38292 5652 38344 5661
rect 3516 5516 3568 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 38292 5176 38344 5228
rect 2228 5108 2280 5160
rect 20 5040 72 5092
rect 4712 4972 4764 5024
rect 36912 5015 36964 5024
rect 36912 4981 36921 5015
rect 36921 4981 36955 5015
rect 36955 4981 36964 5015
rect 36912 4972 36964 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 2688 4632 2740 4684
rect 37096 4675 37148 4684
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 37096 4641 37105 4675
rect 37105 4641 37139 4675
rect 37139 4641 37148 4675
rect 37096 4632 37148 4641
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 25872 4564 25924 4616
rect 38200 4607 38252 4616
rect 38200 4573 38209 4607
rect 38209 4573 38243 4607
rect 38243 4573 38252 4607
rect 38200 4564 38252 4573
rect 3332 4496 3384 4548
rect 19340 4496 19392 4548
rect 38016 4539 38068 4548
rect 38016 4505 38025 4539
rect 38025 4505 38059 4539
rect 38059 4505 38068 4539
rect 38016 4496 38068 4505
rect 3792 4428 3844 4480
rect 5724 4428 5776 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3792 4199 3844 4208
rect 3792 4165 3801 4199
rect 3801 4165 3835 4199
rect 3835 4165 3844 4199
rect 3792 4156 3844 4165
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 24952 4131 25004 4140
rect 24952 4097 24961 4131
rect 24961 4097 24995 4131
rect 24995 4097 25004 4131
rect 24952 4088 25004 4097
rect 37464 4131 37516 4140
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 3148 4020 3200 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8484 4020 8536 4072
rect 2320 3952 2372 4004
rect 37464 4097 37473 4131
rect 37473 4097 37507 4131
rect 37507 4097 37516 4131
rect 37464 4088 37516 4097
rect 35808 4063 35860 4072
rect 35808 4029 35817 4063
rect 35817 4029 35851 4063
rect 35851 4029 35860 4063
rect 35808 4020 35860 4029
rect 4620 3884 4672 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 19432 3884 19484 3936
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 22008 3927 22060 3936
rect 22008 3893 22017 3927
rect 22017 3893 22051 3927
rect 22051 3893 22060 3927
rect 22008 3884 22060 3893
rect 24860 3927 24912 3936
rect 24860 3893 24869 3927
rect 24869 3893 24903 3927
rect 24903 3893 24912 3927
rect 24860 3884 24912 3893
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 30012 3927 30064 3936
rect 30012 3893 30021 3927
rect 30021 3893 30055 3927
rect 30055 3893 30064 3927
rect 30012 3884 30064 3893
rect 33968 3927 34020 3936
rect 33968 3893 33977 3927
rect 33977 3893 34011 3927
rect 34011 3893 34020 3927
rect 33968 3884 34020 3893
rect 34796 3884 34848 3936
rect 37464 3884 37516 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3884 3680 3936 3732
rect 5448 3680 5500 3732
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 3976 3544 4028 3596
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 5632 3612 5684 3664
rect 10876 3612 10928 3664
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 20720 3587 20772 3596
rect 20720 3553 20729 3587
rect 20729 3553 20763 3587
rect 20763 3553 20772 3587
rect 20720 3544 20772 3553
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 25872 3587 25924 3596
rect 25872 3553 25881 3587
rect 25881 3553 25915 3587
rect 25915 3553 25924 3587
rect 25872 3544 25924 3553
rect 26056 3587 26108 3596
rect 26056 3553 26065 3587
rect 26065 3553 26099 3587
rect 26099 3553 26108 3587
rect 26056 3544 26108 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 8852 3476 8904 3528
rect 9772 3476 9824 3528
rect 12900 3476 12952 3528
rect 19340 3476 19392 3528
rect 19984 3476 20036 3528
rect 24308 3476 24360 3528
rect 24584 3476 24636 3528
rect 28264 3476 28316 3528
rect 37372 3612 37424 3664
rect 29092 3544 29144 3596
rect 30012 3587 30064 3596
rect 30012 3553 30021 3587
rect 30021 3553 30055 3587
rect 30055 3553 30064 3587
rect 30012 3544 30064 3553
rect 36268 3544 36320 3596
rect 33876 3519 33928 3528
rect 33876 3485 33885 3519
rect 33885 3485 33919 3519
rect 33919 3485 33928 3519
rect 33876 3476 33928 3485
rect 34796 3476 34848 3528
rect 3240 3451 3292 3460
rect 3240 3417 3249 3451
rect 3249 3417 3283 3451
rect 3283 3417 3292 3451
rect 3240 3408 3292 3417
rect 20904 3451 20956 3460
rect 4344 3340 4396 3392
rect 9036 3340 9088 3392
rect 19340 3340 19392 3392
rect 19524 3340 19576 3392
rect 20904 3417 20913 3451
rect 20913 3417 20947 3451
rect 20947 3417 20956 3451
rect 20904 3408 20956 3417
rect 34060 3408 34112 3460
rect 38660 3408 38712 3460
rect 24400 3340 24452 3392
rect 28080 3340 28132 3392
rect 34152 3340 34204 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 664 3136 716 3188
rect 3516 3111 3568 3120
rect 3516 3077 3525 3111
rect 3525 3077 3559 3111
rect 3559 3077 3568 3111
rect 3516 3068 3568 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 4712 2932 4764 2984
rect 3332 2864 3384 2916
rect 38016 3136 38068 3188
rect 9036 3111 9088 3120
rect 9036 3077 9045 3111
rect 9045 3077 9079 3111
rect 9079 3077 9088 3111
rect 9036 3068 9088 3077
rect 19984 3068 20036 3120
rect 28080 3111 28132 3120
rect 28080 3077 28089 3111
rect 28089 3077 28123 3111
rect 28123 3077 28132 3111
rect 28080 3068 28132 3077
rect 34152 3111 34204 3120
rect 34152 3077 34161 3111
rect 34161 3077 34195 3111
rect 34195 3077 34204 3111
rect 34152 3068 34204 3077
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 11888 3000 11940 3052
rect 12900 3043 12952 3052
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 7472 2932 7524 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 19432 3000 19484 3052
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 33968 3043 34020 3052
rect 33968 3009 33977 3043
rect 33977 3009 34011 3043
rect 34011 3009 34020 3043
rect 33968 3000 34020 3009
rect 36268 3043 36320 3052
rect 36268 3009 36277 3043
rect 36277 3009 36311 3043
rect 36311 3009 36320 3043
rect 36268 3000 36320 3009
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37464 3000 37516 3009
rect 38200 3000 38252 3052
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 22192 2975 22244 2984
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 24492 2975 24544 2984
rect 24492 2941 24501 2975
rect 24501 2941 24535 2975
rect 24535 2941 24544 2975
rect 24492 2932 24544 2941
rect 27896 2975 27948 2984
rect 22008 2864 22060 2916
rect 23204 2864 23256 2916
rect 27896 2941 27905 2975
rect 27905 2941 27939 2975
rect 27939 2941 27948 2975
rect 27896 2932 27948 2941
rect 28356 2975 28408 2984
rect 28356 2941 28365 2975
rect 28365 2941 28399 2975
rect 28399 2941 28408 2975
rect 28356 2932 28408 2941
rect 34796 2975 34848 2984
rect 34796 2941 34805 2975
rect 34805 2941 34839 2975
rect 34839 2941 34848 2975
rect 34796 2932 34848 2941
rect 2596 2796 2648 2848
rect 4712 2796 4764 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3240 2592 3292 2644
rect 6552 2592 6604 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 8392 2592 8444 2644
rect 14740 2592 14792 2644
rect 20904 2592 20956 2644
rect 22192 2592 22244 2644
rect 24492 2592 24544 2644
rect 27896 2592 27948 2644
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2504 2388 2556 2440
rect 4804 2524 4856 2576
rect 4620 2456 4672 2508
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 4712 2456 4764 2465
rect 10876 2524 10928 2576
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 14004 2524 14056 2576
rect 17500 2456 17552 2508
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 24860 2456 24912 2508
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 29920 2456 29972 2508
rect 37188 2524 37240 2576
rect 36912 2499 36964 2508
rect 36912 2465 36921 2499
rect 36921 2465 36955 2499
rect 36955 2465 36964 2499
rect 36912 2456 36964 2465
rect 37648 2456 37700 2508
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 9036 2320 9088 2372
rect 20812 2388 20864 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 29000 2388 29052 2440
rect 17408 2320 17460 2372
rect 28264 2320 28316 2372
rect 30932 2320 30984 2372
rect 9680 2252 9732 2304
rect 17224 2252 17276 2304
rect 17500 2252 17552 2304
rect 24952 2252 25004 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 39200 102 39800
rect 634 39200 746 39800
rect 1278 39200 1390 39800
rect 1922 39200 2034 39800
rect 2566 39200 2678 39800
rect 3210 39200 3322 39800
rect 3854 39200 3966 39800
rect 4498 39200 4610 39800
rect 5142 39200 5254 39800
rect 5786 39200 5898 39800
rect 7074 39200 7186 39800
rect 7718 39200 7830 39800
rect 8362 39200 8474 39800
rect 9006 39200 9118 39800
rect 9650 39200 9762 39800
rect 10294 39200 10406 39800
rect 10938 39200 11050 39800
rect 11582 39200 11694 39800
rect 12226 39200 12338 39800
rect 12452 39222 12756 39250
rect 32 37262 60 39200
rect 1858 37496 1914 37505
rect 1858 37431 1914 37440
rect 20 37256 72 37262
rect 20 37198 72 37204
rect 1872 36854 1900 37431
rect 2412 37324 2464 37330
rect 2412 37266 2464 37272
rect 1860 36848 1912 36854
rect 1860 36790 1912 36796
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1596 35698 1624 36110
rect 1768 36100 1820 36106
rect 1768 36042 1820 36048
rect 1780 35834 1808 36042
rect 1768 35828 1820 35834
rect 1768 35770 1820 35776
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 2424 34610 2452 37266
rect 2504 37256 2556 37262
rect 2504 37198 2556 37204
rect 2516 36854 2544 37198
rect 2504 36848 2556 36854
rect 2504 36790 2556 36796
rect 2608 35894 2636 39200
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2792 36242 2820 38111
rect 3252 36650 3280 39200
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3240 36644 3292 36650
rect 3240 36586 3292 36592
rect 3436 36242 3464 37198
rect 3516 36712 3568 36718
rect 3516 36654 3568 36660
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 3424 36236 3476 36242
rect 3424 36178 3476 36184
rect 2608 35866 2728 35894
rect 2596 35692 2648 35698
rect 2596 35634 2648 35640
rect 2608 34746 2636 35634
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 2412 34604 2464 34610
rect 2412 34546 2464 34552
rect 1860 33992 1912 33998
rect 1860 33934 1912 33940
rect 1872 33522 1900 33934
rect 2044 33856 2096 33862
rect 2044 33798 2096 33804
rect 2056 33590 2084 33798
rect 2044 33584 2096 33590
rect 2044 33526 2096 33532
rect 1860 33516 1912 33522
rect 1860 33458 1912 33464
rect 2504 32496 2556 32502
rect 2504 32438 2556 32444
rect 2516 31822 2544 32438
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 2504 31816 2556 31822
rect 2504 31758 2556 31764
rect 1596 30802 1624 31758
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 30802 1808 31622
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 1584 30796 1636 30802
rect 1584 30738 1636 30744
rect 1768 30796 1820 30802
rect 1768 30738 1820 30744
rect 2136 30048 2188 30054
rect 2136 29990 2188 29996
rect 1584 29572 1636 29578
rect 1584 29514 1636 29520
rect 1596 29345 1624 29514
rect 1582 29336 1638 29345
rect 1582 29271 1638 29280
rect 2148 29170 2176 29990
rect 2136 29164 2188 29170
rect 2136 29106 2188 29112
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1872 28082 1900 28494
rect 1860 28076 1912 28082
rect 1860 28018 1912 28024
rect 2044 28008 2096 28014
rect 2044 27950 2096 27956
rect 2056 27674 2084 27950
rect 2044 27668 2096 27674
rect 2044 27610 2096 27616
rect 1860 22568 1912 22574
rect 1858 22536 1860 22545
rect 1912 22536 1914 22545
rect 1858 22471 1914 22480
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21554 1624 21966
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1596 21010 1624 21111
rect 1584 21004 1636 21010
rect 1584 20946 1636 20952
rect 1952 20528 2004 20534
rect 1950 20496 1952 20505
rect 2004 20496 2006 20505
rect 1950 20431 2006 20440
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1872 17882 1900 18158
rect 2056 17882 2084 18158
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 1860 17128 1912 17134
rect 1858 17096 1860 17105
rect 2136 17128 2188 17134
rect 1912 17096 1914 17105
rect 2136 17070 2188 17076
rect 1858 17031 1914 17040
rect 2148 16794 2176 17070
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2240 16114 2268 18566
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2240 15638 2268 16050
rect 2228 15632 2280 15638
rect 2228 15574 2280 15580
rect 2332 15366 2360 31282
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 2424 23118 2452 27406
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2412 21956 2464 21962
rect 2412 21898 2464 21904
rect 2424 21690 2452 21898
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2516 18834 2544 31758
rect 2608 26234 2636 34682
rect 2700 32366 2728 35866
rect 3528 35834 3556 36654
rect 3896 36258 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4160 37256 4212 37262
rect 4160 37198 4212 37204
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 4172 36786 4200 37198
rect 5356 37188 5408 37194
rect 5356 37130 5408 37136
rect 4344 37120 4396 37126
rect 4344 37062 4396 37068
rect 4356 36854 4384 37062
rect 4344 36848 4396 36854
rect 4344 36790 4396 36796
rect 4160 36780 4212 36786
rect 4160 36722 4212 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3896 36242 4200 36258
rect 3896 36236 4212 36242
rect 3896 36230 4160 36236
rect 4160 36178 4212 36184
rect 4160 36100 4212 36106
rect 4160 36042 4212 36048
rect 4172 35834 4200 36042
rect 3516 35828 3568 35834
rect 3516 35770 3568 35776
rect 4160 35828 4212 35834
rect 4160 35770 4212 35776
rect 3332 35692 3384 35698
rect 3332 35634 3384 35640
rect 3792 35692 3844 35698
rect 3792 35634 3844 35640
rect 3148 34604 3200 34610
rect 3148 34546 3200 34552
rect 2780 33448 2832 33454
rect 2778 33416 2780 33425
rect 2832 33416 2834 33425
rect 2778 33351 2834 33360
rect 2688 32360 2740 32366
rect 2688 32302 2740 32308
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 2780 30796 2832 30802
rect 2780 30738 2832 30744
rect 2792 30705 2820 30738
rect 2778 30696 2834 30705
rect 2778 30631 2834 30640
rect 2872 30592 2924 30598
rect 2872 30534 2924 30540
rect 2884 30054 2912 30534
rect 2872 30048 2924 30054
rect 2872 29990 2924 29996
rect 2884 29594 2912 29990
rect 2976 29714 3004 31078
rect 3160 30258 3188 34546
rect 3344 34542 3372 35634
rect 3332 34536 3384 34542
rect 3332 34478 3384 34484
rect 3240 31204 3292 31210
rect 3240 31146 3292 31152
rect 3148 30252 3200 30258
rect 3148 30194 3200 30200
rect 3056 30116 3108 30122
rect 3056 30058 3108 30064
rect 3068 30025 3096 30058
rect 3054 30016 3110 30025
rect 3054 29951 3110 29960
rect 3160 29866 3188 30194
rect 3068 29838 3188 29866
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 2884 29566 3004 29594
rect 2976 29510 3004 29566
rect 2964 29504 3016 29510
rect 2964 29446 3016 29452
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2872 29096 2924 29102
rect 2872 29038 2924 29044
rect 2792 28762 2820 29038
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2884 28665 2912 29038
rect 2870 28656 2926 28665
rect 2870 28591 2926 28600
rect 2976 28558 3004 29446
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2780 28008 2832 28014
rect 2778 27976 2780 27985
rect 2832 27976 2834 27985
rect 2778 27911 2834 27920
rect 2608 26206 2728 26234
rect 2596 23112 2648 23118
rect 2596 23054 2648 23060
rect 2608 21434 2636 23054
rect 2700 21554 2728 26206
rect 2780 22092 2832 22098
rect 3068 22094 3096 29838
rect 3252 29578 3280 31146
rect 3240 29572 3292 29578
rect 3240 29514 3292 29520
rect 3344 26234 3372 34478
rect 3804 33998 3832 35634
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 3792 33992 3844 33998
rect 3792 33934 3844 33940
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3712 31482 3740 32302
rect 3700 31476 3752 31482
rect 3700 31418 3752 31424
rect 3608 31340 3660 31346
rect 3608 31282 3660 31288
rect 3620 30938 3648 31282
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3620 27470 3648 30874
rect 3608 27464 3660 27470
rect 3608 27406 3660 27412
rect 2780 22034 2832 22040
rect 2976 22066 3096 22094
rect 3160 26206 3372 26234
rect 2792 21865 2820 22034
rect 2778 21856 2834 21865
rect 2778 21791 2834 21800
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2792 21434 2820 21490
rect 2608 21406 2820 21434
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2608 16574 2636 21406
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2700 20058 2728 20334
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2976 18698 3004 22066
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 3068 19990 3096 20810
rect 3056 19984 3108 19990
rect 3056 19926 3108 19932
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2792 17785 2820 18158
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2608 16546 2728 16574
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 1872 14618 1900 14894
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 2240 14074 2268 14894
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2332 12850 2360 13874
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12306 1808 12582
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11762 1624 12174
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9110 2084 9318
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1582 8936 1638 8945
rect 1582 8871 1584 8880
rect 1636 8871 1638 8880
rect 1584 8842 1636 8848
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 8265 1624 8366
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1582 6896 1638 6905
rect 1582 6831 1584 6840
rect 1636 6831 1638 6840
rect 1584 6802 1636 6808
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1872 5234 1900 5646
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 20 5092 72 5098
rect 20 5034 72 5040
rect 32 800 60 5034
rect 2240 4826 2268 5102
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2332 4010 2360 12786
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2424 6458 2452 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 664 3188 716 3194
rect 664 3130 716 3136
rect 676 800 704 3130
rect 1688 2446 1716 3431
rect 2516 2446 2544 6258
rect 2700 4690 2728 16546
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2884 14385 2912 15506
rect 2870 14376 2926 14385
rect 2870 14311 2926 14320
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2778 12336 2834 12345
rect 2778 12271 2780 12280
rect 2832 12271 2834 12280
rect 2780 12242 2832 12248
rect 2884 9586 2912 14214
rect 2976 10674 3004 16390
rect 3068 14414 3096 19382
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3160 13938 3188 26206
rect 3700 23112 3752 23118
rect 3700 23054 3752 23060
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3528 22710 3556 22918
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3712 22642 3740 23054
rect 3700 22636 3752 22642
rect 3700 22578 3752 22584
rect 3804 22094 3832 33934
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3884 32904 3936 32910
rect 3884 32846 3936 32852
rect 3896 32434 3924 32846
rect 3884 32428 3936 32434
rect 3884 32370 3936 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4804 31952 4856 31958
rect 4804 31894 4856 31900
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30258 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30252 4120 30258
rect 4068 30194 4120 30200
rect 4620 30184 4672 30190
rect 4620 30126 4672 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29850 4660 30126
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4632 29034 4660 29582
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4252 28552 4304 28558
rect 4252 28494 4304 28500
rect 4264 28082 4292 28494
rect 4252 28076 4304 28082
rect 4252 28018 4304 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 26784 4028 26790
rect 3976 26726 4028 26732
rect 3988 26450 4016 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4066 26616 4122 26625
rect 4214 26619 4522 26628
rect 4066 26551 4122 26560
rect 4080 26518 4108 26551
rect 4068 26512 4120 26518
rect 4068 26454 4120 26460
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 4160 26308 4212 26314
rect 4160 26250 4212 26256
rect 4172 25786 4200 26250
rect 4080 25758 4200 25786
rect 4080 25498 4108 25758
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 3884 25288 3936 25294
rect 3884 25230 3936 25236
rect 3896 24206 3924 25230
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 4080 24410 4108 24686
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3896 23866 3924 24142
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3712 22066 3832 22094
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3252 21010 3280 21286
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 3620 19310 3648 21422
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3344 18698 3372 18770
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3252 17338 3280 17614
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3252 16182 3280 17274
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3252 14618 3280 15370
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 1676 2440 1728 2446
rect 2504 2440 2556 2446
rect 1676 2382 1728 2388
rect 1858 2408 1914 2417
rect 2504 2382 2556 2388
rect 1858 2343 1860 2352
rect 1912 2343 1914 2352
rect 1860 2314 1912 2320
rect 2608 800 2636 2790
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 2792 785 2820 3538
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2884 1465 2912 2926
rect 2976 2145 3004 4014
rect 3068 2825 3096 11154
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 10810 3280 11018
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9042 3280 9318
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3160 4078 3188 5646
rect 3344 4554 3372 18634
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17270 3556 17478
rect 3516 17264 3568 17270
rect 3516 17206 3568 17212
rect 3620 12434 3648 17682
rect 3712 16182 3740 22066
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3804 20058 3832 20334
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3896 19446 3924 23802
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19848 4120 19854
rect 4066 19816 4068 19825
rect 4120 19816 4122 19825
rect 4066 19751 4122 19760
rect 3884 19440 3936 19446
rect 3884 19382 3936 19388
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3804 16794 3832 19246
rect 3988 18698 4016 19314
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3988 18290 4016 18634
rect 4632 18358 4660 28970
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4724 28626 4752 28902
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 4816 24682 4844 31894
rect 5368 29850 5396 37130
rect 6564 36786 6592 37198
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 7116 36718 7144 39200
rect 9220 37256 9272 37262
rect 9220 37198 9272 37204
rect 9232 36786 9260 37198
rect 9220 36780 9272 36786
rect 9220 36722 9272 36728
rect 9692 36718 9720 39200
rect 6460 36712 6512 36718
rect 6460 36654 6512 36660
rect 7104 36712 7156 36718
rect 7104 36654 7156 36660
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 6472 36378 6500 36654
rect 9416 36378 9444 36654
rect 6460 36372 6512 36378
rect 6460 36314 6512 36320
rect 9404 36372 9456 36378
rect 9404 36314 9456 36320
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6380 35698 6408 36110
rect 8484 36032 8536 36038
rect 8484 35974 8536 35980
rect 6368 35692 6420 35698
rect 6368 35634 6420 35640
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 5356 29844 5408 29850
rect 5356 29786 5408 29792
rect 5368 29170 5396 29786
rect 7668 29646 7696 29990
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7852 28626 7880 28902
rect 5632 28620 5684 28626
rect 5632 28562 5684 28568
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3988 17678 4016 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4724 17678 4752 19722
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4816 17746 4844 18770
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 3988 12434 4016 16730
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 16114 4476 16526
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4540 15348 4568 15642
rect 4632 15502 4660 16050
rect 4724 15706 4752 17614
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4540 15320 4660 15348
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 4080 12714 4108 12951
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3620 12406 3740 12434
rect 3988 12406 4108 12434
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10606 3464 11086
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 6866 3464 7142
rect 3712 6914 3740 12406
rect 3620 6886 3740 6914
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3620 5710 3648 6886
rect 4080 6322 4108 12406
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 3252 2650 3280 3402
rect 3528 3126 3556 5510
rect 4632 5250 4660 15320
rect 4724 9518 4752 15370
rect 4816 15366 4844 16458
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 8974 4752 9454
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4816 6914 4844 15302
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 4724 6886 4844 6914
rect 4724 6390 4752 6886
rect 5368 6866 5396 7142
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4632 5222 4844 5250
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4214 3832 4422
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2962 2136 3018 2145
rect 2962 2071 3018 2080
rect 3344 1714 3372 2858
rect 3252 1686 3372 1714
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 800 3280 1686
rect 3896 800 3924 3674
rect 3988 3602 4016 4558
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 3058 4200 3470
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 3126 4384 3334
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2514 4660 3878
rect 4724 2990 4752 4966
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4724 2514 4752 2790
rect 4816 2582 4844 5222
rect 5460 3738 5488 24686
rect 5644 19854 5672 28562
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 20534 8340 20878
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 8496 16454 8524 35974
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 8944 32360 8996 32366
rect 8944 32302 8996 32308
rect 8956 31890 8984 32302
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 8944 31884 8996 31890
rect 8944 31826 8996 31832
rect 8576 31272 8628 31278
rect 8576 31214 8628 31220
rect 8588 30258 8616 31214
rect 8956 31210 8984 31826
rect 9416 31754 9444 32234
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9956 32224 10008 32230
rect 9956 32166 10008 32172
rect 9404 31748 9456 31754
rect 9404 31690 9456 31696
rect 9312 31680 9364 31686
rect 9312 31622 9364 31628
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 8944 31204 8996 31210
rect 8944 31146 8996 31152
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8956 30054 8984 31146
rect 9048 31142 9076 31282
rect 9324 31278 9352 31622
rect 9692 31346 9720 32166
rect 9968 31822 9996 32166
rect 10428 32026 10456 32846
rect 10508 32768 10560 32774
rect 10508 32710 10560 32716
rect 10520 32434 10548 32710
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10416 32020 10468 32026
rect 10416 31962 10468 31968
rect 9956 31816 10008 31822
rect 9956 31758 10008 31764
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 9036 31136 9088 31142
rect 9036 31078 9088 31084
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 8668 29164 8720 29170
rect 8668 29106 8720 29112
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 8588 26314 8616 26930
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8588 24206 8616 24550
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8680 22098 8708 29106
rect 8760 28416 8812 28422
rect 8760 28358 8812 28364
rect 8772 28014 8800 28358
rect 8852 28076 8904 28082
rect 8852 28018 8904 28024
rect 8760 28008 8812 28014
rect 8760 27950 8812 27956
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8772 25974 8800 26522
rect 8864 26042 8892 28018
rect 8956 26994 8984 29990
rect 9048 29578 9076 31078
rect 9324 30802 9352 31214
rect 9496 31136 9548 31142
rect 9496 31078 9548 31084
rect 9312 30796 9364 30802
rect 9312 30738 9364 30744
rect 9508 30190 9536 31078
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 9588 30320 9640 30326
rect 9588 30262 9640 30268
rect 9496 30184 9548 30190
rect 9496 30126 9548 30132
rect 9404 30116 9456 30122
rect 9404 30058 9456 30064
rect 9128 29776 9180 29782
rect 9128 29718 9180 29724
rect 9036 29572 9088 29578
rect 9036 29514 9088 29520
rect 9140 28558 9168 29718
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9416 27470 9444 30058
rect 9600 29646 9628 30262
rect 10152 30258 10180 30670
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 8956 26382 8984 26930
rect 9232 26586 9260 26930
rect 9312 26920 9364 26926
rect 9312 26862 9364 26868
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 9128 26308 9180 26314
rect 9128 26250 9180 26256
rect 8852 26036 8904 26042
rect 8852 25978 8904 25984
rect 8760 25968 8812 25974
rect 8760 25910 8812 25916
rect 9140 24070 9168 26250
rect 9324 25906 9352 26862
rect 9404 26784 9456 26790
rect 9404 26726 9456 26732
rect 9416 26450 9444 26726
rect 9600 26586 9628 27474
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9404 26444 9456 26450
rect 9404 26386 9456 26392
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9600 25906 9628 26318
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 9416 24410 9444 24822
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9048 23730 9076 24006
rect 9140 23730 9168 24006
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8680 21554 8708 22034
rect 8864 21554 8892 23462
rect 9048 23118 9076 23666
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9600 22574 9628 23054
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9692 22094 9720 29038
rect 9772 24880 9824 24886
rect 9772 24822 9824 24828
rect 9784 23730 9812 24822
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9692 22066 9812 22094
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 8680 21010 8708 21490
rect 8668 21004 8720 21010
rect 8668 20946 8720 20952
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8588 20466 8616 20742
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8680 20262 8708 20946
rect 8864 20942 8892 21490
rect 9140 21146 9168 21490
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8864 20602 8892 20878
rect 9600 20874 9628 21422
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9692 20874 9720 21286
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9600 20754 9628 20810
rect 9600 20726 9720 20754
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8864 18290 8892 18770
rect 9140 18766 9168 20266
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9140 18290 9168 18702
rect 9324 18698 9628 18714
rect 9324 18692 9640 18698
rect 9324 18686 9588 18692
rect 9324 18630 9352 18686
rect 9588 18634 9640 18640
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9600 18290 9628 18634
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 8864 17678 8892 18226
rect 9140 17882 9168 18226
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8864 16590 8892 17614
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 6458 5580 6666
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5552 3602 5580 3878
rect 5644 3670 5672 15914
rect 9140 13802 9168 16594
rect 9600 15502 9628 18226
rect 9692 18222 9720 20726
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 17746 9720 18158
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9784 17252 9812 22066
rect 9876 19242 9904 22442
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9876 18970 9904 19178
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17678 9904 18022
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9968 17252 9996 30126
rect 10152 29714 10180 30194
rect 10140 29708 10192 29714
rect 10140 29650 10192 29656
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10060 29306 10088 29582
rect 10048 29300 10100 29306
rect 10048 29242 10100 29248
rect 10152 29170 10180 29650
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10232 24200 10284 24206
rect 10284 24160 10364 24188
rect 10232 24142 10284 24148
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 10060 23798 10088 24074
rect 10048 23792 10100 23798
rect 10048 23734 10100 23740
rect 10060 23202 10088 23734
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 10152 23322 10180 23666
rect 10336 23526 10364 24160
rect 10428 24138 10456 24550
rect 10416 24132 10468 24138
rect 10416 24074 10468 24080
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10060 23174 10180 23202
rect 10336 23186 10364 23462
rect 10152 23118 10180 23174
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10060 21962 10088 22918
rect 10612 22681 10640 32846
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 12176 32026 12204 32302
rect 12164 32020 12216 32026
rect 12164 31962 12216 31968
rect 11796 31884 11848 31890
rect 11796 31826 11848 31832
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11072 30734 11100 31214
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10980 29170 11008 29786
rect 10968 29164 11020 29170
rect 10968 29106 11020 29112
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 11072 27538 11100 27882
rect 11164 27606 11192 28018
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10796 26586 10824 27406
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10796 26382 10824 26522
rect 10888 26382 10916 26726
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 11072 26042 11100 26250
rect 11716 26234 11744 31214
rect 11808 29170 11836 31826
rect 12452 31754 12480 39222
rect 12728 39114 12756 39222
rect 12870 39200 12982 39800
rect 14158 39200 14270 39800
rect 14802 39200 14914 39800
rect 15446 39200 15558 39800
rect 16090 39200 16202 39800
rect 16734 39200 16846 39800
rect 17378 39200 17490 39800
rect 18022 39200 18134 39800
rect 18666 39200 18778 39800
rect 19310 39200 19422 39800
rect 19954 39200 20066 39800
rect 20598 39200 20710 39800
rect 21886 39200 21998 39800
rect 22530 39200 22642 39800
rect 23174 39200 23286 39800
rect 23818 39200 23930 39800
rect 24462 39200 24574 39800
rect 25106 39200 25218 39800
rect 25750 39200 25862 39800
rect 26394 39200 26506 39800
rect 27038 39200 27150 39800
rect 27682 39200 27794 39800
rect 28970 39200 29082 39800
rect 29614 39200 29726 39800
rect 30258 39200 30370 39800
rect 30902 39200 31014 39800
rect 31546 39200 31658 39800
rect 32190 39200 32302 39800
rect 32834 39200 32946 39800
rect 33478 39200 33590 39800
rect 34122 39200 34234 39800
rect 34766 39200 34878 39800
rect 35410 39200 35522 39800
rect 36698 39200 36810 39800
rect 37342 39200 37454 39800
rect 37986 39200 38098 39800
rect 38630 39200 38742 39800
rect 39274 39200 39386 39800
rect 12912 39114 12940 39200
rect 12728 39086 12940 39114
rect 14464 37256 14516 37262
rect 14464 37198 14516 37204
rect 14476 36242 14504 37198
rect 14648 37120 14700 37126
rect 14648 37062 14700 37068
rect 14660 36854 14688 37062
rect 14648 36848 14700 36854
rect 14648 36790 14700 36796
rect 14464 36236 14516 36242
rect 14464 36178 14516 36184
rect 14648 35012 14700 35018
rect 14648 34954 14700 34960
rect 14464 34400 14516 34406
rect 14464 34342 14516 34348
rect 14476 33998 14504 34342
rect 14660 34202 14688 34954
rect 14844 34746 14872 39200
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 14936 36718 14964 37198
rect 14924 36712 14976 36718
rect 14924 36654 14976 36660
rect 16132 36242 16160 39200
rect 16212 37256 16264 37262
rect 16212 37198 16264 37204
rect 16120 36236 16172 36242
rect 16120 36178 16172 36184
rect 14924 36100 14976 36106
rect 14924 36042 14976 36048
rect 14936 35834 14964 36042
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15212 35834 15240 35974
rect 16224 35894 16252 37198
rect 16776 36854 16804 39200
rect 16764 36848 16816 36854
rect 16764 36790 16816 36796
rect 17420 36242 17448 39200
rect 17592 37256 17644 37262
rect 17592 37198 17644 37204
rect 17604 36922 17632 37198
rect 17592 36916 17644 36922
rect 17592 36858 17644 36864
rect 18064 36718 18092 39200
rect 19156 37324 19208 37330
rect 19156 37266 19208 37272
rect 18880 37256 18932 37262
rect 18880 37198 18932 37204
rect 18696 37120 18748 37126
rect 18696 37062 18748 37068
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 18708 36242 18736 37062
rect 18892 36242 18920 37198
rect 19168 36786 19196 37266
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19444 36786 19472 37198
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 20640 36718 20668 39200
rect 21928 37618 21956 39200
rect 22572 38026 22600 39200
rect 22572 37998 22876 38026
rect 21928 37590 22048 37618
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 18972 36712 19024 36718
rect 18972 36654 19024 36660
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 20628 36712 20680 36718
rect 20628 36654 20680 36660
rect 17408 36236 17460 36242
rect 17408 36178 17460 36184
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 18880 36236 18932 36242
rect 18880 36178 18932 36184
rect 16224 35866 16344 35894
rect 14924 35828 14976 35834
rect 14924 35770 14976 35776
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 15212 35698 15240 35770
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 15292 35624 15344 35630
rect 15292 35566 15344 35572
rect 15304 35086 15332 35566
rect 15384 35216 15436 35222
rect 15384 35158 15436 35164
rect 15292 35080 15344 35086
rect 15292 35022 15344 35028
rect 14832 34740 14884 34746
rect 14832 34682 14884 34688
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 14740 34468 14792 34474
rect 14740 34410 14792 34416
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14752 33454 14780 34410
rect 15120 33930 15148 34478
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 15120 33522 15148 33866
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 14740 33448 14792 33454
rect 14740 33390 14792 33396
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 12716 32768 12768 32774
rect 12716 32710 12768 32716
rect 12728 32434 12756 32710
rect 12716 32428 12768 32434
rect 12716 32370 12768 32376
rect 13544 32224 13596 32230
rect 13544 32166 13596 32172
rect 13556 31754 13584 32166
rect 13912 31952 13964 31958
rect 13912 31894 13964 31900
rect 12452 31726 12572 31754
rect 11980 30252 12032 30258
rect 12164 30252 12216 30258
rect 11980 30194 12032 30200
rect 12084 30212 12164 30240
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11900 29306 11928 29990
rect 11992 29850 12020 30194
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 11992 29578 12020 29786
rect 11980 29572 12032 29578
rect 11980 29514 12032 29520
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11808 28762 11836 29106
rect 11888 28960 11940 28966
rect 11888 28902 11940 28908
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 11900 28626 11928 28902
rect 11888 28620 11940 28626
rect 11888 28562 11940 28568
rect 11992 28558 12020 29514
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 11980 28416 12032 28422
rect 12084 28370 12112 30212
rect 12164 30194 12216 30200
rect 12164 30116 12216 30122
rect 12164 30058 12216 30064
rect 12176 29102 12204 30058
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 12452 29306 12480 29582
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12164 29096 12216 29102
rect 12164 29038 12216 29044
rect 12176 28762 12204 29038
rect 12164 28756 12216 28762
rect 12164 28698 12216 28704
rect 12032 28364 12112 28370
rect 11980 28358 12112 28364
rect 11992 28342 12112 28358
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11808 27674 11836 27950
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11992 26790 12020 28342
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11992 26382 12020 26726
rect 12176 26382 12204 28698
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12360 26790 12388 26930
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 11716 26206 11928 26234
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11808 24410 11836 25842
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10704 23118 10732 24074
rect 11808 23798 11836 24346
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 10876 23588 10928 23594
rect 10876 23530 10928 23536
rect 10888 23118 10916 23530
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10598 22672 10654 22681
rect 10598 22607 10654 22616
rect 10704 22030 10732 23054
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10704 20874 10732 21966
rect 10692 20868 10744 20874
rect 10692 20810 10744 20816
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10244 19378 10272 19654
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18970 10180 19110
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10152 18834 10180 18906
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10244 18766 10272 19314
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10336 18970 10364 19246
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 9692 17224 9812 17252
rect 9876 17224 9996 17252
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 12850 9168 13738
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9508 12986 9536 13194
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5736 3602 5764 4422
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 5828 800 5856 6802
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4162 8340 4558
rect 8220 4146 8340 4162
rect 8208 4140 8340 4146
rect 8260 4134 8340 4140
rect 8208 4082 8260 4088
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6564 2650 6592 2926
rect 7484 2650 7512 2926
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7760 800 7788 2926
rect 8404 2650 8432 4014
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8496 2258 8524 4014
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8864 3058 8892 3470
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 3126 9076 3334
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 8404 2230 8524 2258
rect 8404 800 8432 2230
rect 9048 800 9076 2314
rect 9692 2310 9720 17224
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9784 11762 9812 15302
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9876 6914 9904 17224
rect 10244 16590 10272 18702
rect 10336 18290 10364 18906
rect 10692 18896 10744 18902
rect 10690 18864 10692 18873
rect 10744 18864 10746 18873
rect 10690 18799 10746 18808
rect 10796 18766 10824 19246
rect 11072 18766 11100 19382
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10796 17678 10824 18702
rect 11164 18426 11192 19246
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 16114 10272 16526
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10244 14074 10272 14282
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10060 13530 10088 13874
rect 10336 13530 10364 15506
rect 10428 14414 10456 17614
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10520 16046 10548 16594
rect 11808 16522 11836 18226
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10520 15910 10548 15982
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 11440 15706 11468 16390
rect 11808 16046 11836 16458
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11532 15706 11560 15914
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10336 12986 10364 13466
rect 10428 13394 10456 14350
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9968 11218 9996 12650
rect 10244 12306 10272 12786
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10336 12238 10364 12922
rect 10428 12850 10456 13194
rect 10704 12918 10732 13194
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 11256 12782 11284 13262
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10520 12442 10548 12582
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11286 10548 11698
rect 11808 11626 11836 12174
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9784 6886 9904 6914
rect 9784 3534 9812 6886
rect 10520 4146 10548 11222
rect 11624 11218 11652 11494
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 10612 3602 10640 3878
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10888 2582 10916 3606
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10980 800 11008 3538
rect 11808 2514 11836 3878
rect 11900 3058 11928 26206
rect 12452 25906 12480 29242
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12544 24274 12572 31726
rect 13544 31748 13596 31754
rect 13544 31690 13596 31696
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 13084 30252 13136 30258
rect 13084 30194 13136 30200
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 12636 26450 12664 26930
rect 12728 26858 12756 29446
rect 13096 27538 13124 30194
rect 13372 29578 13400 30670
rect 13556 30258 13584 31690
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13740 30326 13768 30534
rect 13728 30320 13780 30326
rect 13728 30262 13780 30268
rect 13544 30252 13596 30258
rect 13544 30194 13596 30200
rect 13924 30122 13952 31894
rect 14200 31482 14228 32846
rect 14648 32836 14700 32842
rect 14648 32778 14700 32784
rect 14660 32570 14688 32778
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14188 31476 14240 31482
rect 14188 31418 14240 31424
rect 14292 30938 14320 31758
rect 14752 31142 14780 33390
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14844 32434 14872 33254
rect 14924 32768 14976 32774
rect 14924 32710 14976 32716
rect 14832 32428 14884 32434
rect 14832 32370 14884 32376
rect 14936 31958 14964 32710
rect 15028 32434 15056 33458
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 15120 32230 15148 33458
rect 15304 32994 15332 35022
rect 15396 34610 15424 35158
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 15384 34604 15436 34610
rect 15384 34546 15436 34552
rect 15672 34066 15700 34886
rect 15936 34740 15988 34746
rect 15936 34682 15988 34688
rect 15660 34060 15712 34066
rect 15660 34002 15712 34008
rect 15212 32966 15332 32994
rect 15212 32910 15240 32966
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 14924 31952 14976 31958
rect 14924 31894 14976 31900
rect 15120 31346 15148 32166
rect 15212 31890 15240 32846
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15108 31340 15160 31346
rect 15108 31282 15160 31288
rect 14740 31136 14792 31142
rect 14740 31078 14792 31084
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 14280 30932 14332 30938
rect 14280 30874 14332 30880
rect 15028 30802 15056 31078
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 15016 30796 15068 30802
rect 15016 30738 15068 30744
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13648 29646 13676 29990
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 13360 29572 13412 29578
rect 13360 29514 13412 29520
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13820 29504 13872 29510
rect 13820 29446 13872 29452
rect 13280 28082 13308 29446
rect 13832 29102 13860 29446
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13924 28966 13952 30058
rect 14292 29782 14320 30738
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14280 29776 14332 29782
rect 14280 29718 14332 29724
rect 14476 29646 14504 30194
rect 15120 30054 15148 31282
rect 15212 30802 15240 31826
rect 15672 31686 15700 34002
rect 15384 31680 15436 31686
rect 15384 31622 15436 31628
rect 15660 31680 15712 31686
rect 15660 31622 15712 31628
rect 15292 31204 15344 31210
rect 15292 31146 15344 31152
rect 15304 30870 15332 31146
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 15304 30648 15332 30806
rect 15212 30620 15332 30648
rect 15212 30394 15240 30620
rect 15200 30388 15252 30394
rect 15200 30330 15252 30336
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 15108 30048 15160 30054
rect 15108 29990 15160 29996
rect 14936 29646 14964 29990
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 14292 29102 14320 29582
rect 14752 29102 14780 29582
rect 15120 29170 15148 29990
rect 15292 29776 15344 29782
rect 15292 29718 15344 29724
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 15304 29034 15332 29718
rect 15396 29646 15424 31622
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15856 30938 15884 31282
rect 15844 30932 15896 30938
rect 15844 30874 15896 30880
rect 15856 30394 15884 30874
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15672 29714 15700 30262
rect 15856 30122 15884 30330
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 15396 28966 15424 29582
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15580 29034 15608 29446
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15476 29028 15528 29034
rect 15476 28970 15528 28976
rect 15568 29028 15620 29034
rect 15568 28970 15620 28976
rect 13912 28960 13964 28966
rect 13912 28902 13964 28908
rect 15384 28960 15436 28966
rect 15384 28902 15436 28908
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 13372 27606 13400 27950
rect 13360 27600 13412 27606
rect 13360 27542 13412 27548
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 15396 27470 15424 28018
rect 15488 27470 15516 28970
rect 15580 28014 15608 28970
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15672 27470 15700 29038
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15764 27878 15792 28970
rect 15948 28234 15976 34682
rect 16028 32428 16080 32434
rect 16028 32370 16080 32376
rect 16040 31890 16068 32370
rect 16028 31884 16080 31890
rect 16028 31826 16080 31832
rect 16040 31346 16068 31826
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 16040 30326 16068 31282
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 15948 28206 16068 28234
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15764 27470 15792 27814
rect 13912 27464 13964 27470
rect 13912 27406 13964 27412
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15660 27464 15712 27470
rect 15660 27406 15712 27412
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12716 26852 12768 26858
rect 12716 26794 12768 26800
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12728 26042 12756 26794
rect 12820 26586 12848 26930
rect 13924 26926 13952 27406
rect 15672 27334 15700 27406
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 12900 26240 12952 26246
rect 12900 26182 12952 26188
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12728 25498 12756 25842
rect 12716 25492 12768 25498
rect 12716 25434 12768 25440
rect 12912 25294 12940 26182
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13740 24410 13768 24686
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12268 23118 12296 23734
rect 12360 23730 12388 24142
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13372 23730 13400 24006
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12360 23050 12388 23666
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 13464 22642 13492 23462
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13740 22778 13768 23190
rect 13832 23118 13860 23802
rect 13924 23662 13952 26862
rect 14280 26376 14332 26382
rect 15672 26364 15700 27270
rect 15936 26444 15988 26450
rect 15936 26386 15988 26392
rect 15844 26376 15896 26382
rect 15672 26336 15844 26364
rect 14280 26318 14332 26324
rect 15844 26318 15896 26324
rect 14292 26042 14320 26318
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14292 25770 14320 25978
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 14280 25764 14332 25770
rect 14280 25706 14332 25712
rect 14924 25764 14976 25770
rect 14924 25706 14976 25712
rect 14936 25498 14964 25706
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 15212 25294 15240 25774
rect 15764 25498 15792 26182
rect 15948 26042 15976 26386
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15752 25492 15804 25498
rect 15752 25434 15804 25440
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14108 23866 14136 24142
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14292 23730 14320 24346
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 12452 21894 12480 22578
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22030 12756 22510
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12992 21956 13044 21962
rect 12992 21898 13044 21904
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12452 21622 12480 21830
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11992 19854 12020 21490
rect 13004 21486 13032 21898
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11992 18970 12020 19790
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 12176 18358 12204 20878
rect 12360 18426 12388 21286
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 20602 12480 20810
rect 13004 20806 13032 21422
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 13096 20262 13124 22170
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13188 21350 13216 21966
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13188 21146 13216 21286
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13188 20534 13216 21082
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13280 20466 13308 21286
rect 13464 21010 13492 21966
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13464 20466 13492 20946
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12452 16590 12480 18226
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 16726 12664 17206
rect 13004 17202 13032 18022
rect 13096 17882 13124 20198
rect 13464 19514 13492 20402
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13464 19258 13492 19450
rect 13464 19230 13584 19258
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13464 18970 13492 19110
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13556 18766 13584 19230
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13648 18902 13676 19110
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13740 18086 13768 22714
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 21418 13860 21490
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13924 20466 13952 23598
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 14108 21554 14136 22170
rect 14200 22098 14228 23598
rect 14292 23254 14320 23666
rect 14384 23322 14412 24686
rect 15212 24070 15240 25230
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15476 23792 15528 23798
rect 15476 23734 15528 23740
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14280 23248 14332 23254
rect 14280 23190 14332 23196
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14752 22098 14780 22918
rect 15488 22778 15516 23734
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14200 21418 14228 22034
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14384 21554 14412 21898
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14384 20942 14412 21490
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 20942 14504 21422
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 14476 19854 14504 20878
rect 14660 20262 14688 20946
rect 14844 20262 14872 22578
rect 15488 22234 15516 22714
rect 15672 22642 15700 23666
rect 15856 23322 15884 25842
rect 15936 25356 15988 25362
rect 15936 25298 15988 25304
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15028 22030 15056 22170
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 14936 21486 14964 21966
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15120 21554 15148 21830
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15488 21486 15516 22170
rect 15672 22098 15700 22578
rect 15856 22438 15884 23258
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15580 21690 15608 21898
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 15212 19854 15240 21354
rect 15856 21350 15884 22374
rect 15948 21554 15976 25298
rect 16040 24818 16068 28206
rect 16212 28144 16264 28150
rect 16212 28086 16264 28092
rect 16224 27674 16252 28086
rect 16212 27668 16264 27674
rect 16212 27610 16264 27616
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16132 25838 16160 26386
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 16132 23118 16160 24006
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16132 22710 16160 23054
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15856 19786 15884 21286
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 14464 19712 14516 19718
rect 14462 19680 14464 19689
rect 14516 19680 14518 19689
rect 14462 19615 14518 19624
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 12912 16794 12940 17002
rect 13188 16794 13216 17002
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 13556 16590 13584 17206
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 16794 13676 17138
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 12452 16250 12480 16526
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 15026 12480 15302
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12532 14952 12584 14958
rect 12636 14940 12664 16458
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 14958 12756 15846
rect 12584 14912 12664 14940
rect 12532 14894 12584 14900
rect 12636 14074 12664 14912
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12820 14822 12848 16186
rect 13372 15162 13400 16526
rect 13740 15502 13768 18022
rect 13832 17678 13860 18702
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14568 17882 14596 18634
rect 15028 18222 15056 19178
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 15028 17678 15056 18158
rect 15212 17678 15240 18566
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 13832 17202 13860 17614
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14200 16658 14228 16934
rect 14476 16794 14504 16934
rect 14660 16794 14688 17138
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14936 16046 14964 17478
rect 15304 16998 15332 19382
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 18290 15792 18566
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15856 18154 15884 19722
rect 15948 19718 15976 21490
rect 16316 20058 16344 35866
rect 18984 35834 19012 36654
rect 19904 36378 19932 36654
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 21008 36242 21036 37198
rect 20996 36236 21048 36242
rect 22020 36224 22048 37590
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22284 37120 22336 37126
rect 22284 37062 22336 37068
rect 22296 36854 22324 37062
rect 22284 36848 22336 36854
rect 22284 36790 22336 36796
rect 22756 36718 22784 37198
rect 22848 36718 22876 37998
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 22744 36712 22796 36718
rect 22744 36654 22796 36660
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22100 36236 22152 36242
rect 22020 36196 22100 36224
rect 20996 36178 21048 36184
rect 22100 36178 22152 36184
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 18972 35828 19024 35834
rect 18972 35770 19024 35776
rect 16948 35692 17000 35698
rect 16948 35634 17000 35640
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 16960 35290 16988 35634
rect 17868 35488 17920 35494
rect 17868 35430 17920 35436
rect 16948 35284 17000 35290
rect 16948 35226 17000 35232
rect 17592 35080 17644 35086
rect 17592 35022 17644 35028
rect 17604 34746 17632 35022
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17880 34542 17908 35430
rect 18892 35290 18920 35634
rect 18696 35284 18748 35290
rect 18696 35226 18748 35232
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18144 34944 18196 34950
rect 18144 34886 18196 34892
rect 18156 34610 18184 34886
rect 18420 34672 18472 34678
rect 18420 34614 18472 34620
rect 18144 34604 18196 34610
rect 18144 34546 18196 34552
rect 17408 34536 17460 34542
rect 17408 34478 17460 34484
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 16856 33992 16908 33998
rect 16856 33934 16908 33940
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16592 32842 16620 33798
rect 16868 33658 16896 33934
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 16580 32836 16632 32842
rect 16580 32778 16632 32784
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16684 30326 16712 31758
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16776 29306 16804 32778
rect 17420 32434 17448 34478
rect 18156 34202 18184 34546
rect 18432 34202 18460 34614
rect 18708 34406 18736 35226
rect 18788 35012 18840 35018
rect 18788 34954 18840 34960
rect 18880 35012 18932 35018
rect 18880 34954 18932 34960
rect 18696 34400 18748 34406
rect 18696 34342 18748 34348
rect 18144 34196 18196 34202
rect 18144 34138 18196 34144
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 17972 33590 18000 33934
rect 17960 33584 18012 33590
rect 17960 33526 18012 33532
rect 18156 33522 18184 34138
rect 18708 33998 18736 34342
rect 18800 33998 18828 34954
rect 18892 34678 18920 34954
rect 19352 34746 19380 36110
rect 21180 36100 21232 36106
rect 21180 36042 21232 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 21192 35834 21220 36042
rect 23296 36032 23348 36038
rect 23296 35974 23348 35980
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 23308 35766 23336 35974
rect 23296 35760 23348 35766
rect 23296 35702 23348 35708
rect 23492 35698 23520 36858
rect 23584 36786 23612 37198
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23860 36650 23888 39200
rect 23848 36644 23900 36650
rect 23848 36586 23900 36592
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 23480 35692 23532 35698
rect 23480 35634 23532 35640
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 18880 34672 18932 34678
rect 18880 34614 18932 34620
rect 18696 33992 18748 33998
rect 18696 33934 18748 33940
rect 18788 33992 18840 33998
rect 18788 33934 18840 33940
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18708 33810 18736 33934
rect 18892 33862 18920 34614
rect 18972 34536 19024 34542
rect 18972 34478 19024 34484
rect 18880 33856 18932 33862
rect 18144 33516 18196 33522
rect 18144 33458 18196 33464
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17604 32434 17632 32710
rect 17408 32428 17460 32434
rect 17408 32370 17460 32376
rect 17592 32428 17644 32434
rect 17592 32370 17644 32376
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17236 30938 17264 31214
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17328 30734 17356 32166
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 17328 30394 17356 30670
rect 17408 30660 17460 30666
rect 17408 30602 17460 30608
rect 17420 30394 17448 30602
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16868 27962 16896 29514
rect 16960 29458 16988 29990
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 16960 29430 17080 29458
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 16960 29102 16988 29242
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16960 28762 16988 29038
rect 16948 28756 17000 28762
rect 16948 28698 17000 28704
rect 16776 27934 16896 27962
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16684 24138 16712 25094
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16500 23322 16528 23462
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16776 20806 16804 27934
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27062 16896 27814
rect 16856 27056 16908 27062
rect 16856 26998 16908 27004
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23866 16988 24006
rect 16948 23860 17000 23866
rect 16948 23802 17000 23808
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16868 20618 16896 22578
rect 16776 20602 16896 20618
rect 16960 20602 16988 23802
rect 17052 22982 17080 29430
rect 17144 29170 17172 29582
rect 17236 29306 17264 30126
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 17144 25362 17172 29106
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17236 26042 17264 26794
rect 17328 26790 17356 28562
rect 17420 28558 17448 30330
rect 17604 30122 17632 31758
rect 18064 31278 18092 33390
rect 18524 32434 18552 33798
rect 18708 33782 18828 33810
rect 18880 33798 18932 33804
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18616 32842 18644 33526
rect 18800 32910 18828 33782
rect 18984 33454 19012 34478
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19260 33658 19288 33934
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 18972 33448 19024 33454
rect 18972 33390 19024 33396
rect 18788 32904 18840 32910
rect 18788 32846 18840 32852
rect 18604 32836 18656 32842
rect 18604 32778 18656 32784
rect 18696 32836 18748 32842
rect 18696 32778 18748 32784
rect 18616 32434 18644 32778
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18604 32428 18656 32434
rect 18604 32370 18656 32376
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18144 31748 18196 31754
rect 18144 31690 18196 31696
rect 18156 31482 18184 31690
rect 18144 31476 18196 31482
rect 18144 31418 18196 31424
rect 18340 31278 18368 31758
rect 18420 31680 18472 31686
rect 18420 31622 18472 31628
rect 18432 31346 18460 31622
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18340 30734 18368 31214
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 17972 30326 18000 30670
rect 18236 30592 18288 30598
rect 18236 30534 18288 30540
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 17500 30116 17552 30122
rect 17500 30058 17552 30064
rect 17592 30116 17644 30122
rect 17592 30058 17644 30064
rect 17512 29782 17540 30058
rect 17500 29776 17552 29782
rect 17972 29730 18000 30262
rect 17500 29718 17552 29724
rect 17788 29702 18000 29730
rect 17788 29646 17816 29702
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 17132 25220 17184 25226
rect 17132 25162 17184 25168
rect 17144 23186 17172 25162
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16764 20596 16896 20602
rect 16816 20590 16896 20596
rect 16948 20596 17000 20602
rect 16764 20538 16816 20544
rect 16948 20538 17000 20544
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16856 19984 16908 19990
rect 16856 19926 16908 19932
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 16040 17898 16068 19314
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16132 18290 16160 18362
rect 16316 18290 16344 18702
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16040 17870 16160 17898
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16590 15332 16934
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14936 15570 14964 15982
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13556 15026 13584 15370
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12636 13802 12664 14010
rect 12728 13938 12756 14214
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11762 12020 12038
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12268 11354 12296 13262
rect 12544 12306 12572 13398
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12360 11354 12388 12242
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12544 11830 12572 12106
rect 12636 12102 12664 13738
rect 12728 12782 12756 13874
rect 12820 13462 12848 14758
rect 13280 13530 13308 14962
rect 13556 13938 13584 14962
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14346 14136 14758
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 14200 14074 14228 14962
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 13280 12646 13308 13466
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12728 12238 12756 12582
rect 13372 12442 13400 13262
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12986 14228 13194
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13464 12442 13492 12650
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12912 11898 12940 12242
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12622 11384 12678 11393
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12348 11348 12400 11354
rect 12622 11319 12624 11328
rect 12348 11290 12400 11296
rect 12676 11319 12678 11328
rect 12624 11290 12676 11296
rect 12728 11150 12756 11494
rect 12912 11354 12940 11834
rect 14016 11762 14044 12786
rect 14200 12374 14228 12922
rect 14292 12918 14320 14214
rect 14660 14074 14688 14826
rect 14936 14414 14964 15506
rect 15488 15502 15516 15846
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14660 13938 14688 14010
rect 15580 13938 15608 17750
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16040 16590 16068 17138
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 16114 15700 16390
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 16132 14890 16160 17870
rect 16212 17808 16264 17814
rect 16212 17750 16264 17756
rect 16224 16998 16252 17750
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 15502 16252 16934
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16132 14482 16160 14826
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13938 16160 14214
rect 16224 14074 16252 14282
rect 16316 14074 16344 14350
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 14648 13932 14700 13938
rect 14568 13892 14648 13920
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14568 12714 14596 13892
rect 14648 13874 14700 13880
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13530 14780 13806
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14200 11898 14228 12310
rect 14660 12238 14688 12854
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15304 12714 15332 12786
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14660 11762 14688 12174
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12912 3058 12940 3470
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12268 800 12296 2450
rect 13556 800 13584 2926
rect 14016 2582 14044 11698
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14476 11150 14504 11562
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14752 2650 14780 12174
rect 15580 11762 15608 12310
rect 15672 12306 15700 12786
rect 16132 12782 16160 13874
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 12306 15792 12582
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15764 11830 15792 12242
rect 16224 12238 16252 12650
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16132 11898 16160 12174
rect 16224 12102 16252 12174
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 15856 11354 15884 11698
rect 16224 11558 16252 11698
rect 16408 11626 16436 19858
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16592 17610 16620 18294
rect 16684 18290 16712 19654
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 13870 16528 15302
rect 16684 14618 16712 17682
rect 16776 16794 16804 18158
rect 16868 17542 16896 19926
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16960 17270 16988 19246
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 17052 17066 17080 20742
rect 17144 20262 17172 21286
rect 17236 20942 17264 21558
rect 17224 20936 17276 20942
rect 17222 20904 17224 20913
rect 17276 20904 17278 20913
rect 17222 20839 17278 20848
rect 17328 20754 17356 26726
rect 17420 26586 17448 26998
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17408 26240 17460 26246
rect 17408 26182 17460 26188
rect 17420 25702 17448 26182
rect 17604 25974 17632 26318
rect 17592 25968 17644 25974
rect 17592 25910 17644 25916
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 24206 17540 24550
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17604 23866 17632 24074
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17696 23594 17724 27882
rect 18144 27396 18196 27402
rect 18144 27338 18196 27344
rect 18156 27130 18184 27338
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 18064 25498 18092 25910
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 18248 25294 18276 30534
rect 18340 30326 18368 30670
rect 18328 30320 18380 30326
rect 18328 30262 18380 30268
rect 18616 29714 18644 32370
rect 18708 30802 18736 32778
rect 18800 32230 18828 32846
rect 19444 32434 19472 35022
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34610 20024 34886
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 20076 34536 20128 34542
rect 20128 34484 20208 34490
rect 20076 34478 20208 34484
rect 20088 34462 20208 34478
rect 20180 34406 20208 34462
rect 20168 34400 20220 34406
rect 20168 34342 20220 34348
rect 20180 34202 20208 34342
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 19904 33425 19932 33458
rect 19890 33416 19946 33425
rect 19890 33351 19946 33360
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19996 32910 20024 33254
rect 20088 33046 20116 33458
rect 20076 33040 20128 33046
rect 20076 32982 20128 32988
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19996 32366 20024 32710
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 19984 32360 20036 32366
rect 19984 32302 20036 32308
rect 18788 32224 18840 32230
rect 19168 32212 19196 32302
rect 19616 32224 19668 32230
rect 19168 32184 19288 32212
rect 18788 32166 18840 32172
rect 18696 30796 18748 30802
rect 18696 30738 18748 30744
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18604 29708 18656 29714
rect 18604 29650 18656 29656
rect 18708 29238 18736 30534
rect 18800 29578 18828 32166
rect 19260 31634 19288 32184
rect 19616 32166 19668 32172
rect 19628 32026 19656 32166
rect 19616 32020 19668 32026
rect 19616 31962 19668 31968
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19812 31822 19840 31962
rect 19800 31816 19852 31822
rect 19800 31758 19852 31764
rect 20088 31754 20116 32982
rect 20076 31748 20128 31754
rect 20076 31690 20128 31696
rect 19340 31680 19392 31686
rect 19260 31628 19340 31634
rect 19260 31622 19392 31628
rect 19260 31606 19380 31622
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 18788 29572 18840 29578
rect 18788 29514 18840 29520
rect 18800 29238 18828 29514
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 18788 29232 18840 29238
rect 18788 29174 18840 29180
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 19076 28914 19104 30738
rect 19156 30184 19208 30190
rect 19156 30126 19208 30132
rect 19168 29034 19196 30126
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 18432 27538 18460 28902
rect 19076 28886 19196 28914
rect 19168 28490 19196 28886
rect 19156 28484 19208 28490
rect 19156 28426 19208 28432
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 17776 25288 17828 25294
rect 18236 25288 18288 25294
rect 17776 25230 17828 25236
rect 18064 25248 18236 25276
rect 17684 23588 17736 23594
rect 17684 23530 17736 23536
rect 17788 23118 17816 25230
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17592 22704 17644 22710
rect 17592 22646 17644 22652
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17420 22098 17448 22578
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17420 21146 17448 22034
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17236 20726 17356 20754
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17144 19922 17172 20198
rect 17126 19916 17178 19922
rect 17126 19858 17178 19864
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17144 19514 17172 19654
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17236 19446 17264 20726
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18970 17264 19246
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17328 18834 17356 20198
rect 17420 19854 17448 20538
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17144 18290 17172 18566
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16868 16250 16896 16594
rect 16960 16590 16988 16934
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17052 15434 17080 16050
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16500 12918 16528 13806
rect 16684 13802 16712 14554
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16684 13462 16712 13738
rect 16960 13530 16988 13874
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 17144 13326 17172 18090
rect 17236 16250 17264 18294
rect 17328 18154 17356 18566
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17328 17270 17356 17682
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17420 16794 17448 18566
rect 17512 17626 17540 21830
rect 17604 20942 17632 22646
rect 17696 22094 17724 22918
rect 17788 22778 17816 23054
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 17880 22710 17908 22986
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17868 22094 17920 22098
rect 17696 22092 17920 22094
rect 17696 22066 17868 22092
rect 17868 22034 17920 22040
rect 17972 21622 18000 24754
rect 18064 23118 18092 25248
rect 18236 25230 18288 25236
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18156 23798 18184 24006
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 18156 23662 18184 23693
rect 18144 23656 18196 23662
rect 18340 23610 18368 26794
rect 19168 26518 19196 28426
rect 19260 26994 19288 31606
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19352 30258 19380 30670
rect 19444 30326 19472 31078
rect 20088 30734 20116 31690
rect 20076 30728 20128 30734
rect 20076 30670 20128 30676
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19800 30320 19852 30326
rect 19800 30262 19852 30268
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19444 29594 19472 30262
rect 19708 30048 19760 30054
rect 19812 30002 19840 30262
rect 20088 30258 20116 30670
rect 20076 30252 20128 30258
rect 20076 30194 20128 30200
rect 19892 30116 19944 30122
rect 19892 30058 19944 30064
rect 19760 29996 19840 30002
rect 19708 29990 19840 29996
rect 19720 29974 19840 29990
rect 19812 29850 19840 29974
rect 19800 29844 19852 29850
rect 19800 29786 19852 29792
rect 19904 29646 19932 30058
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19892 29640 19944 29646
rect 19444 29578 19564 29594
rect 19892 29582 19944 29588
rect 19444 29572 19576 29578
rect 19444 29566 19524 29572
rect 19524 29514 19576 29520
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19444 27538 19472 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19892 28212 19944 28218
rect 19892 28154 19944 28160
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19444 27334 19472 27474
rect 19628 27470 19656 27814
rect 19904 27674 19932 28154
rect 19996 27946 20024 29990
rect 20088 29646 20116 30194
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 20076 29504 20128 29510
rect 20076 29446 20128 29452
rect 20088 28014 20116 29446
rect 20180 28778 20208 34138
rect 20442 33416 20498 33425
rect 20260 33380 20312 33386
rect 20442 33351 20498 33360
rect 20260 33322 20312 33328
rect 20272 32892 20300 33322
rect 20352 32904 20404 32910
rect 20272 32864 20352 32892
rect 20272 32366 20300 32864
rect 20352 32846 20404 32852
rect 20260 32360 20312 32366
rect 20260 32302 20312 32308
rect 20272 31890 20300 32302
rect 20260 31884 20312 31890
rect 20260 31826 20312 31832
rect 20456 30802 20484 33351
rect 20628 33312 20680 33318
rect 20628 33254 20680 33260
rect 20536 32292 20588 32298
rect 20536 32234 20588 32240
rect 20548 31890 20576 32234
rect 20640 32026 20668 33254
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20640 31890 20668 31962
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20548 31142 20576 31690
rect 20732 31414 20760 35634
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 21272 35080 21324 35086
rect 21272 35022 21324 35028
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 21008 34746 21036 35022
rect 20996 34740 21048 34746
rect 20996 34682 21048 34688
rect 21284 34082 21312 35022
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22388 34678 22416 34886
rect 22376 34672 22428 34678
rect 22376 34614 22428 34620
rect 21284 34054 21496 34082
rect 21468 33998 21496 34054
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 22388 33946 22416 34614
rect 22928 34604 22980 34610
rect 22928 34546 22980 34552
rect 22468 33992 22520 33998
rect 22388 33940 22468 33946
rect 22388 33934 22520 33940
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 21272 33924 21324 33930
rect 21272 33866 21324 33872
rect 21008 33114 21036 33866
rect 21088 33856 21140 33862
rect 21088 33798 21140 33804
rect 21100 33522 21128 33798
rect 21284 33658 21312 33866
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 21272 33448 21324 33454
rect 21178 33416 21234 33425
rect 21272 33390 21324 33396
rect 21178 33351 21234 33360
rect 20996 33108 21048 33114
rect 20996 33050 21048 33056
rect 21192 32910 21220 33351
rect 21284 32978 21312 33390
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21376 33046 21404 33254
rect 21364 33040 21416 33046
rect 21364 32982 21416 32988
rect 21272 32972 21324 32978
rect 21272 32914 21324 32920
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21364 32904 21416 32910
rect 21364 32846 21416 32852
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 20824 31822 20852 32370
rect 21376 32366 21404 32846
rect 21364 32360 21416 32366
rect 21364 32302 21416 32308
rect 21468 31890 21496 33934
rect 22388 33918 22508 33934
rect 22388 32910 22416 33918
rect 22836 33856 22888 33862
rect 22836 33798 22888 33804
rect 22848 32910 22876 33798
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 22468 32836 22520 32842
rect 22468 32778 22520 32784
rect 22480 32366 22508 32778
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22480 31958 22508 32302
rect 22468 31952 22520 31958
rect 22468 31894 22520 31900
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 20812 31816 20864 31822
rect 20864 31764 20944 31770
rect 20812 31758 20944 31764
rect 20824 31742 20944 31758
rect 20720 31408 20772 31414
rect 20720 31350 20772 31356
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20628 30864 20680 30870
rect 20628 30806 20680 30812
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20456 29646 20484 30738
rect 20640 29850 20668 30806
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20916 29646 20944 31742
rect 21008 31754 21036 31826
rect 21008 31726 21128 31754
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 20180 28750 20392 28778
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 20180 28082 20208 28426
rect 20272 28150 20300 28630
rect 20260 28144 20312 28150
rect 20260 28086 20312 28092
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20076 28008 20128 28014
rect 20076 27950 20128 27956
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19156 26512 19208 26518
rect 19156 26454 19208 26460
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18616 25770 18644 26318
rect 18604 25764 18656 25770
rect 18604 25706 18656 25712
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18420 25220 18472 25226
rect 18420 25162 18472 25168
rect 18432 24818 18460 25162
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18524 24206 18552 25298
rect 18616 25294 18644 25706
rect 19168 25362 19196 26454
rect 19156 25356 19208 25362
rect 19156 25298 19208 25304
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18196 23604 18368 23610
rect 18144 23598 18368 23604
rect 18156 23582 18368 23598
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17604 20466 17632 20878
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17604 18630 17632 20402
rect 17684 19440 17736 19446
rect 17684 19382 17736 19388
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17696 18426 17724 19382
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17604 18086 17632 18226
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17512 17598 17724 17626
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17236 13938 17264 16186
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 17144 12646 17172 13262
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17236 12238 17264 13874
rect 17328 12442 17356 16050
rect 17512 13326 17540 17138
rect 17604 16590 17632 17478
rect 17696 16946 17724 17598
rect 17788 17270 17816 21354
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17972 20534 18000 20742
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 17972 19718 18000 20266
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17866 18864 17922 18873
rect 17866 18799 17922 18808
rect 17880 18698 17908 18799
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17972 16998 18000 19654
rect 18064 19242 18092 23054
rect 18156 20058 18184 23582
rect 18432 23474 18460 23666
rect 18248 23446 18460 23474
rect 18248 22778 18276 23446
rect 18420 23248 18472 23254
rect 18420 23190 18472 23196
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 18432 22438 18460 23190
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18052 19236 18104 19242
rect 18052 19178 18104 19184
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18156 17882 18184 18294
rect 18248 18222 18276 21286
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18340 19514 18368 19722
rect 18432 19530 18460 22374
rect 18512 21956 18564 21962
rect 18512 21898 18564 21904
rect 18524 20942 18552 21898
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18328 19508 18380 19514
rect 18432 19502 18552 19530
rect 18328 19450 18380 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18432 18358 18460 19314
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 17960 16992 18012 16998
rect 17696 16918 17816 16946
rect 17960 16934 18012 16940
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17696 16590 17724 16730
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17604 15366 17632 16526
rect 17696 15502 17724 16526
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17512 12986 17540 13262
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17604 12918 17632 14214
rect 17788 13258 17816 16918
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15638 18000 16050
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 18248 15570 18276 16390
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18432 14618 18460 18294
rect 18524 18154 18552 19502
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18524 17678 18552 18090
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18432 13734 18460 14554
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18524 13530 18552 16526
rect 18616 16182 18644 25230
rect 19352 24410 19380 26862
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19444 25702 19472 26182
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18800 23866 18828 24142
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18800 22982 18828 23802
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 21350 18828 22918
rect 19444 22094 19472 25298
rect 19904 25294 19932 25638
rect 19996 25498 20024 26250
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24206 20116 24754
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19352 22066 19472 22094
rect 19352 21434 19380 22066
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 19260 21406 19380 21434
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 19174 18736 19790
rect 18800 19718 18828 20946
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18984 20466 19012 20742
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19260 20346 19288 21406
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20466 19380 21286
rect 19812 20874 19840 21490
rect 19996 20942 20024 22510
rect 20088 22030 20116 23258
rect 20180 23254 20208 28018
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20272 27470 20300 27882
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20272 27130 20300 27406
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20088 21078 20116 21966
rect 20272 21418 20300 26318
rect 20364 24682 20392 28750
rect 20824 28558 20852 29582
rect 21100 29170 21128 31726
rect 21180 31272 21232 31278
rect 21180 31214 21232 31220
rect 21192 29170 21220 31214
rect 22100 30728 22152 30734
rect 22100 30670 22152 30676
rect 22112 29850 22140 30670
rect 22376 30660 22428 30666
rect 22376 30602 22428 30608
rect 22388 30122 22416 30602
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22376 30116 22428 30122
rect 22376 30058 22428 30064
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 20628 26512 20680 26518
rect 20628 26454 20680 26460
rect 20640 25974 20668 26454
rect 20628 25968 20680 25974
rect 20628 25910 20680 25916
rect 20824 25294 20852 28494
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20916 27402 20944 28358
rect 21008 27470 21036 28494
rect 20996 27464 21048 27470
rect 20996 27406 21048 27412
rect 20904 27396 20956 27402
rect 20904 27338 20956 27344
rect 20916 27282 20944 27338
rect 20916 27254 21036 27282
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20916 25906 20944 26318
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 20732 23866 20760 24754
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20364 21554 20392 22986
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20548 22234 20576 22578
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20640 22094 20668 23530
rect 20718 22672 20774 22681
rect 20718 22607 20720 22616
rect 20772 22607 20774 22616
rect 20720 22578 20772 22584
rect 20732 22234 20760 22578
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20548 22066 20668 22094
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20534 19472 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19996 20398 20024 20878
rect 19984 20392 20036 20398
rect 19260 20318 19380 20346
rect 19984 20334 20036 20340
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18788 19712 18840 19718
rect 18892 19689 18920 19722
rect 18788 19654 18840 19660
rect 18878 19680 18934 19689
rect 18878 19615 18934 19624
rect 19352 19446 19380 20318
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18708 15570 18736 19110
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 19168 15162 19196 17682
rect 19352 17134 19380 19382
rect 19444 17202 19472 19722
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 17678 20024 19654
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 20180 18970 20208 19382
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20364 17814 20392 18702
rect 20352 17808 20404 17814
rect 20352 17750 20404 17756
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19996 17066 20024 17614
rect 20548 17218 20576 22066
rect 20824 20942 20852 24006
rect 20904 23792 20956 23798
rect 20902 23760 20904 23769
rect 20956 23760 20958 23769
rect 20902 23695 20958 23704
rect 21008 22094 21036 27254
rect 21100 23186 21128 29106
rect 21192 29050 21220 29106
rect 21192 29022 21312 29050
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 21192 28558 21220 28902
rect 21284 28626 21312 29022
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21284 27538 21312 28562
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21272 27532 21324 27538
rect 21272 27474 21324 27480
rect 21732 27328 21784 27334
rect 21732 27270 21784 27276
rect 21364 26784 21416 26790
rect 21364 26726 21416 26732
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 20916 22066 21036 22094
rect 20916 22030 20944 22066
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20916 21690 20944 21966
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20916 20754 20944 21626
rect 20824 20726 20944 20754
rect 20824 20602 20852 20726
rect 21192 20618 21220 22170
rect 21284 22030 21312 25094
rect 21376 24614 21404 26726
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21376 21690 21404 22510
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20916 20590 21220 20618
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19854 20760 20198
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 19378 20760 19654
rect 20824 19446 20852 20538
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20824 18970 20852 19246
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20640 18426 20668 18702
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20824 18290 20852 18566
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20364 17190 20576 17218
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 15502 19288 15846
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19168 13938 19196 15098
rect 19260 14006 19288 15438
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15162 20116 15370
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19996 15026 20024 15098
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14414 19472 14758
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14074 20024 14554
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 14074 20116 14214
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13818 19196 13874
rect 19168 13790 19380 13818
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17788 12918 17816 13194
rect 17972 12986 18000 13330
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17420 12374 17448 12786
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17604 12238 17632 12854
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18156 12374 18184 12786
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18248 12238 18276 12786
rect 18432 12442 18460 12786
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 17236 11694 17264 12174
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17328 11694 17356 11834
rect 18432 11694 18460 12174
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 16224 11014 16252 11494
rect 16316 11150 16344 11494
rect 16408 11218 16436 11562
rect 17236 11286 17264 11630
rect 18524 11393 18552 13466
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19260 12850 19288 12922
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19260 12594 19288 12786
rect 19352 12782 19380 13790
rect 19444 12850 19472 14010
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20180 12986 20208 15302
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 19340 12776 19392 12782
rect 19392 12724 19472 12730
rect 19340 12718 19472 12724
rect 19352 12702 19472 12718
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11830 18920 12174
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 19168 11626 19196 12582
rect 19260 12566 19380 12594
rect 19352 12102 19380 12566
rect 19444 12170 19472 12702
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 12442 20024 12582
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11762 19380 12038
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20088 11762 20116 12106
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 18510 11384 18566 11393
rect 18420 11348 18472 11354
rect 18510 11319 18566 11328
rect 18420 11290 18472 11296
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 18340 10674 18368 11018
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18432 10062 18460 11290
rect 18524 11286 18552 11319
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 19812 11218 19840 11698
rect 20180 11558 20208 12786
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20272 11694 20300 12174
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 20180 11150 20208 11494
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 18616 10266 18644 10542
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 3534 19380 4490
rect 19444 4026 19472 10542
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20364 8498 20392 17190
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 12442 20576 14894
rect 20536 12436 20588 12442
rect 20916 12434 20944 20590
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21192 20058 21220 20402
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21008 18358 21036 19790
rect 21468 19514 21496 19790
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21100 18086 21128 18702
rect 21192 18222 21220 19246
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17202 21036 17614
rect 21100 17270 21128 18022
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21192 17202 21220 17682
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21744 16590 21772 27270
rect 21836 26382 21864 28494
rect 22756 28082 22784 30126
rect 22940 28218 22968 34546
rect 23400 34202 23428 35022
rect 24504 34542 24532 39200
rect 24584 36712 24636 36718
rect 24584 36654 24636 36660
rect 24596 36378 24624 36654
rect 24584 36372 24636 36378
rect 24584 36314 24636 36320
rect 25148 36242 25176 39200
rect 25792 37330 25820 39200
rect 25780 37324 25832 37330
rect 26436 37312 26464 39200
rect 26436 37284 26556 37312
rect 25780 37266 25832 37272
rect 26240 37188 26292 37194
rect 26240 37130 26292 37136
rect 26424 37188 26476 37194
rect 26424 37130 26476 37136
rect 26252 36922 26280 37130
rect 26240 36916 26292 36922
rect 26240 36858 26292 36864
rect 25136 36236 25188 36242
rect 25136 36178 25188 36184
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24596 35698 24624 36110
rect 24768 36100 24820 36106
rect 24768 36042 24820 36048
rect 24780 35834 24808 36042
rect 25044 36032 25096 36038
rect 25044 35974 25096 35980
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 25056 35698 25084 35974
rect 26436 35834 26464 37130
rect 26528 36650 26556 37284
rect 26516 36644 26568 36650
rect 26516 36586 26568 36592
rect 27080 36242 27108 39200
rect 27344 36712 27396 36718
rect 27344 36654 27396 36660
rect 27068 36236 27120 36242
rect 27068 36178 27120 36184
rect 26884 36168 26936 36174
rect 26884 36110 26936 36116
rect 26608 36100 26660 36106
rect 26608 36042 26660 36048
rect 26424 35828 26476 35834
rect 26424 35770 26476 35776
rect 24584 35692 24636 35698
rect 24584 35634 24636 35640
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 25964 35692 26016 35698
rect 25964 35634 26016 35640
rect 25056 35154 25084 35634
rect 25044 35148 25096 35154
rect 25044 35090 25096 35096
rect 25976 34950 26004 35634
rect 26620 35290 26648 36042
rect 26896 35290 26924 36110
rect 27356 35766 27384 36654
rect 27724 35766 27752 39200
rect 28632 37324 28684 37330
rect 28632 37266 28684 37272
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 27816 36854 27844 37198
rect 27804 36848 27856 36854
rect 27804 36790 27856 36796
rect 28448 36644 28500 36650
rect 28448 36586 28500 36592
rect 27344 35760 27396 35766
rect 27344 35702 27396 35708
rect 27712 35760 27764 35766
rect 27712 35702 27764 35708
rect 27988 35624 28040 35630
rect 27988 35566 28040 35572
rect 28000 35290 28028 35566
rect 26608 35284 26660 35290
rect 26608 35226 26660 35232
rect 26884 35284 26936 35290
rect 26884 35226 26936 35232
rect 27988 35284 28040 35290
rect 27988 35226 28040 35232
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 25412 34944 25464 34950
rect 25412 34886 25464 34892
rect 25964 34944 26016 34950
rect 25964 34886 26016 34892
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23768 33658 23796 34478
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 23756 33652 23808 33658
rect 23756 33594 23808 33600
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 23664 33516 23716 33522
rect 23664 33458 23716 33464
rect 23676 33386 23704 33458
rect 23664 33380 23716 33386
rect 23664 33322 23716 33328
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 23124 30326 23152 30534
rect 23388 30388 23440 30394
rect 23388 30330 23440 30336
rect 23112 30320 23164 30326
rect 23112 30262 23164 30268
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23032 29714 23060 30194
rect 23020 29708 23072 29714
rect 23020 29650 23072 29656
rect 23400 29170 23428 30330
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 23492 29578 23520 30194
rect 23480 29572 23532 29578
rect 23480 29514 23532 29520
rect 23388 29164 23440 29170
rect 23388 29106 23440 29112
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 22928 28212 22980 28218
rect 22928 28154 22980 28160
rect 23216 28082 23244 28358
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 22756 27062 22784 28018
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 23032 27470 23060 27814
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22744 27056 22796 27062
rect 22744 26998 22796 27004
rect 22756 26586 22784 26998
rect 22940 26790 22968 27270
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 22744 26580 22796 26586
rect 22744 26522 22796 26528
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21836 25770 21864 26318
rect 23400 25906 23428 29106
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23492 26994 23520 27814
rect 23572 27396 23624 27402
rect 23572 27338 23624 27344
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23584 26382 23612 27338
rect 23676 26874 23704 33322
rect 24504 32570 24532 33526
rect 24584 33312 24636 33318
rect 24584 33254 24636 33260
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24412 31346 24440 31622
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 23756 29572 23808 29578
rect 23756 29514 23808 29520
rect 23768 28150 23796 29514
rect 24044 29238 24072 30194
rect 24032 29232 24084 29238
rect 24032 29174 24084 29180
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23768 27402 23796 28086
rect 24044 27878 24072 28154
rect 24412 28082 24440 28358
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 24044 27470 24072 27814
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 24032 27328 24084 27334
rect 24032 27270 24084 27276
rect 23860 27062 23888 27270
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 23940 26920 23992 26926
rect 23676 26846 23888 26874
rect 23940 26862 23992 26868
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 21824 25764 21876 25770
rect 21824 25706 21876 25712
rect 21836 25362 21864 25706
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22296 24750 22324 25230
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22296 23798 22324 24686
rect 22480 24410 22508 25162
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22664 24274 22692 25842
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22848 24818 22876 25162
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23216 24954 23244 25094
rect 23204 24948 23256 24954
rect 23204 24890 23256 24896
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22112 23254 22140 23666
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22100 23248 22152 23254
rect 22100 23190 22152 23196
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22778 21956 22918
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22204 22642 22232 23598
rect 22296 23186 22324 23734
rect 22836 23520 22888 23526
rect 22836 23462 22888 23468
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22756 22710 22784 22918
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22204 22094 22232 22578
rect 22112 22066 22232 22094
rect 21914 21448 21970 21457
rect 21914 21383 21916 21392
rect 21968 21383 21970 21392
rect 21916 21354 21968 21360
rect 22112 21078 22140 22066
rect 22100 21072 22152 21078
rect 22020 21020 22100 21026
rect 22020 21014 22152 21020
rect 22020 20998 22140 21014
rect 22020 20466 22048 20998
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22112 17610 22140 20878
rect 22296 20466 22324 22646
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22664 19786 22692 21490
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22204 18766 22232 19722
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22480 18902 22508 19314
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22388 18698 22416 18838
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21008 14822 21036 16390
rect 21284 16114 21312 16390
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21100 14618 21128 14962
rect 21284 14822 21312 15030
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21836 14346 21864 16390
rect 22020 16114 22048 17478
rect 22388 17202 22416 18634
rect 22480 18426 22508 18838
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22756 18426 22784 18770
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21928 13530 21956 15098
rect 22020 14482 22048 16050
rect 22848 14890 22876 23462
rect 23124 17882 23152 24142
rect 23216 24138 23244 24890
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 23216 21622 23244 24074
rect 23584 24070 23612 26318
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23572 23180 23624 23186
rect 23572 23122 23624 23128
rect 23584 22964 23612 23122
rect 23676 23118 23704 24822
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23768 22982 23796 24142
rect 23756 22976 23808 22982
rect 23584 22936 23704 22964
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23400 20942 23428 22374
rect 23584 21486 23612 22442
rect 23676 21894 23704 22936
rect 23756 22918 23808 22924
rect 23768 22030 23796 22918
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23204 20324 23256 20330
rect 23204 20266 23256 20272
rect 23216 19310 23244 20266
rect 23676 19854 23704 21354
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23216 18766 23244 19246
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 23032 17202 23060 17546
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23124 17270 23152 17478
rect 23216 17338 23244 18566
rect 23492 18290 23520 19110
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23584 18086 23612 19654
rect 23676 19310 23704 19790
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23768 19242 23796 21490
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23860 18698 23888 26846
rect 23952 26586 23980 26862
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 23952 23866 23980 26522
rect 24044 26382 24072 27270
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 24320 26382 24348 26726
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24044 25498 24072 26318
rect 24596 25498 24624 33254
rect 24688 32434 24716 33798
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24768 32836 24820 32842
rect 24768 32778 24820 32784
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24688 31346 24716 32370
rect 24780 31686 24808 32778
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24676 31340 24728 31346
rect 24676 31282 24728 31288
rect 24780 30122 24808 31622
rect 24872 31414 24900 31962
rect 24964 31482 24992 32914
rect 25136 32836 25188 32842
rect 25136 32778 25188 32784
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 24860 31408 24912 31414
rect 24860 31350 24912 31356
rect 24768 30116 24820 30122
rect 24768 30058 24820 30064
rect 24872 29850 24900 31350
rect 25056 31346 25084 32166
rect 25148 31482 25176 32778
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25320 32360 25372 32366
rect 25320 32302 25372 32308
rect 25240 31958 25268 32302
rect 25332 32026 25360 32302
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25228 31952 25280 31958
rect 25228 31894 25280 31900
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 25056 30938 25084 31282
rect 25044 30932 25096 30938
rect 25044 30874 25096 30880
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24676 29708 24728 29714
rect 24676 29650 24728 29656
rect 24688 26874 24716 29650
rect 25424 29102 25452 34886
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 25504 33924 25556 33930
rect 25504 33866 25556 33872
rect 25516 33658 25544 33866
rect 25504 33652 25556 33658
rect 25504 33594 25556 33600
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 25608 33046 25636 33526
rect 25596 33040 25648 33046
rect 25596 32982 25648 32988
rect 25504 32292 25556 32298
rect 25504 32234 25556 32240
rect 25516 31822 25544 32234
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 25608 30938 25636 31282
rect 25596 30932 25648 30938
rect 25596 30874 25648 30880
rect 25884 30802 25912 31282
rect 25872 30796 25924 30802
rect 25872 30738 25924 30744
rect 25976 30274 26004 33934
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 26068 32570 26096 32846
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26252 31482 26280 32846
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 26148 31408 26200 31414
rect 26148 31350 26200 31356
rect 26160 30802 26188 31350
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 26252 30666 26280 31282
rect 26528 30938 26556 35022
rect 28460 34474 28488 36586
rect 28644 35766 28672 37266
rect 29012 36242 29040 39200
rect 29656 36802 29684 39200
rect 30300 37330 30328 39200
rect 30288 37324 30340 37330
rect 30288 37266 30340 37272
rect 30104 37188 30156 37194
rect 30104 37130 30156 37136
rect 29656 36774 29776 36802
rect 29748 36718 29776 36774
rect 29644 36712 29696 36718
rect 29644 36654 29696 36660
rect 29736 36712 29788 36718
rect 29736 36654 29788 36660
rect 29000 36236 29052 36242
rect 29000 36178 29052 36184
rect 29092 36168 29144 36174
rect 29092 36110 29144 36116
rect 28632 35760 28684 35766
rect 28632 35702 28684 35708
rect 29104 34474 29132 36110
rect 29656 35290 29684 36654
rect 29920 36100 29972 36106
rect 29920 36042 29972 36048
rect 29932 35834 29960 36042
rect 29920 35828 29972 35834
rect 29920 35770 29972 35776
rect 30116 35290 30144 37130
rect 30656 37120 30708 37126
rect 30656 37062 30708 37068
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 30564 35692 30616 35698
rect 30564 35634 30616 35640
rect 29644 35284 29696 35290
rect 29644 35226 29696 35232
rect 30104 35284 30156 35290
rect 30104 35226 30156 35232
rect 30208 35222 30236 35634
rect 30196 35216 30248 35222
rect 30196 35158 30248 35164
rect 30576 34746 30604 35634
rect 30668 35290 30696 37062
rect 30944 36242 30972 39200
rect 31760 36848 31812 36854
rect 31760 36790 31812 36796
rect 30932 36236 30984 36242
rect 30932 36178 30984 36184
rect 31772 35290 31800 36790
rect 32232 36650 32260 39200
rect 32876 37330 32904 39200
rect 32864 37324 32916 37330
rect 32864 37266 32916 37272
rect 33048 37324 33100 37330
rect 33048 37266 33100 37272
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 32312 36712 32364 36718
rect 32312 36654 32364 36660
rect 32220 36644 32272 36650
rect 32220 36586 32272 36592
rect 32036 36168 32088 36174
rect 32036 36110 32088 36116
rect 32048 35698 32076 36110
rect 32220 36100 32272 36106
rect 32220 36042 32272 36048
rect 32232 35834 32260 36042
rect 32220 35828 32272 35834
rect 32220 35770 32272 35776
rect 32036 35692 32088 35698
rect 32036 35634 32088 35640
rect 32324 35290 32352 36654
rect 30656 35284 30708 35290
rect 30656 35226 30708 35232
rect 31760 35284 31812 35290
rect 31760 35226 31812 35232
rect 32312 35284 32364 35290
rect 32312 35226 32364 35232
rect 32312 35012 32364 35018
rect 32312 34954 32364 34960
rect 30564 34740 30616 34746
rect 30564 34682 30616 34688
rect 28448 34468 28500 34474
rect 28448 34410 28500 34416
rect 29092 34468 29144 34474
rect 29092 34410 29144 34416
rect 26976 34060 27028 34066
rect 26976 34002 27028 34008
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 26804 33454 26832 33934
rect 26988 33522 27016 34002
rect 27252 33992 27304 33998
rect 27252 33934 27304 33940
rect 27896 33992 27948 33998
rect 27896 33934 27948 33940
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 26792 33448 26844 33454
rect 26792 33390 26844 33396
rect 26700 33040 26752 33046
rect 26700 32982 26752 32988
rect 26608 32768 26660 32774
rect 26608 32710 26660 32716
rect 26620 32434 26648 32710
rect 26608 32428 26660 32434
rect 26608 32370 26660 32376
rect 26712 31210 26740 32982
rect 26700 31204 26752 31210
rect 26700 31146 26752 31152
rect 26516 30932 26568 30938
rect 26516 30874 26568 30880
rect 26240 30660 26292 30666
rect 26240 30602 26292 30608
rect 26056 30320 26108 30326
rect 25976 30268 26056 30274
rect 25976 30262 26108 30268
rect 25976 30246 26096 30262
rect 25976 29238 26004 30246
rect 26252 29850 26280 30602
rect 26528 30394 26556 30874
rect 26700 30864 26752 30870
rect 26700 30806 26752 30812
rect 26516 30388 26568 30394
rect 26516 30330 26568 30336
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 26240 29844 26292 29850
rect 26240 29786 26292 29792
rect 26528 29646 26556 30126
rect 26712 29714 26740 30806
rect 26804 30734 26832 33390
rect 26884 32972 26936 32978
rect 26884 32914 26936 32920
rect 26896 32502 26924 32914
rect 26988 32910 27016 33458
rect 27068 33108 27120 33114
rect 27068 33050 27120 33056
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 26884 32496 26936 32502
rect 27080 32450 27108 33050
rect 27172 32774 27200 33798
rect 27264 33658 27292 33934
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27264 32966 27476 32994
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 26884 32438 26936 32444
rect 26988 32422 27108 32450
rect 27172 32434 27200 32710
rect 27264 32434 27292 32966
rect 27448 32910 27476 32966
rect 27908 32910 27936 33934
rect 27988 33516 28040 33522
rect 27988 33458 28040 33464
rect 27344 32904 27396 32910
rect 27344 32846 27396 32852
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 27160 32428 27212 32434
rect 26988 31890 27016 32422
rect 27160 32370 27212 32376
rect 27252 32428 27304 32434
rect 27252 32370 27304 32376
rect 27068 32360 27120 32366
rect 27068 32302 27120 32308
rect 27080 32026 27108 32302
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 26988 31346 27016 31826
rect 27264 31414 27292 32370
rect 27356 32314 27384 32846
rect 27528 32768 27580 32774
rect 27528 32710 27580 32716
rect 27540 32434 27568 32710
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 27356 32286 27568 32314
rect 28000 32298 28028 33458
rect 28172 33312 28224 33318
rect 28172 33254 28224 33260
rect 28184 32978 28212 33254
rect 28172 32972 28224 32978
rect 28172 32914 28224 32920
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 27540 31754 27568 32286
rect 27988 32292 28040 32298
rect 27988 32234 28040 32240
rect 28000 32026 28028 32234
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 27252 31408 27304 31414
rect 27252 31350 27304 31356
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 27344 31204 27396 31210
rect 27344 31146 27396 31152
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 27252 30728 27304 30734
rect 27252 30670 27304 30676
rect 26700 29708 26752 29714
rect 26700 29650 26752 29656
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 25964 29232 26016 29238
rect 25964 29174 26016 29180
rect 25412 29096 25464 29102
rect 25412 29038 25464 29044
rect 26332 29028 26384 29034
rect 26332 28970 26384 28976
rect 25228 28552 25280 28558
rect 25228 28494 25280 28500
rect 25240 27946 25268 28494
rect 25504 28484 25556 28490
rect 25504 28426 25556 28432
rect 25228 27940 25280 27946
rect 25228 27882 25280 27888
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24872 26994 24900 27338
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24688 26846 24808 26874
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 24688 26382 24716 26726
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24032 25492 24084 25498
rect 24032 25434 24084 25440
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24780 25430 24808 26846
rect 24860 26852 24912 26858
rect 24860 26794 24912 26800
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24780 25294 24808 25366
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24872 25140 24900 26794
rect 24964 26314 24992 26930
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24780 25112 24900 25140
rect 24780 24614 24808 25112
rect 24860 24880 24912 24886
rect 24860 24822 24912 24828
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24872 24070 24900 24822
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 23940 23860 23992 23866
rect 23940 23802 23992 23808
rect 23952 22094 23980 23802
rect 24780 23730 24808 24006
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 24872 23186 24900 24006
rect 24964 23798 24992 26250
rect 25240 25770 25268 27882
rect 25516 26858 25544 28426
rect 26344 28422 26372 28970
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 26344 28082 26372 28358
rect 26436 28218 26464 28902
rect 26528 28762 26556 29582
rect 26516 28756 26568 28762
rect 26516 28698 26568 28704
rect 26424 28212 26476 28218
rect 26424 28154 26476 28160
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26528 28014 26556 28698
rect 26516 28008 26568 28014
rect 26516 27950 26568 27956
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25700 27130 25728 27270
rect 25688 27124 25740 27130
rect 25688 27066 25740 27072
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25504 26852 25556 26858
rect 25504 26794 25556 26800
rect 25792 26586 25820 26930
rect 25780 26580 25832 26586
rect 25780 26522 25832 26528
rect 25228 25764 25280 25770
rect 25228 25706 25280 25712
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25148 24274 25176 24550
rect 25516 24410 25544 24550
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 24216 23044 24268 23050
rect 24216 22986 24268 22992
rect 24228 22098 24256 22986
rect 23952 22066 24072 22094
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23952 21554 23980 21830
rect 24044 21690 24072 22066
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24124 21956 24176 21962
rect 24124 21898 24176 21904
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24136 21554 24164 21898
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24044 19854 24072 20334
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 24044 19446 24072 19790
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24136 19378 24164 19722
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 24136 18630 24164 19314
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23676 17338 23704 18226
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 16998 23060 17138
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23216 15638 23244 17274
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23308 16590 23336 17138
rect 23388 17128 23440 17134
rect 23440 17076 23612 17082
rect 23388 17070 23612 17076
rect 23400 17066 23612 17070
rect 23400 17060 23624 17066
rect 23400 17054 23572 17060
rect 23572 17002 23624 17008
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23768 16538 23796 16934
rect 23308 16250 23336 16526
rect 23768 16510 23888 16538
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 23584 15570 23612 15982
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23584 15162 23612 15506
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22020 14006 22048 14418
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 20536 12378 20588 12384
rect 20824 12406 20944 12434
rect 20824 11014 20852 12406
rect 21836 12238 21864 13262
rect 22112 12442 22140 14350
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 13530 22232 14214
rect 22388 13938 22416 14486
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22756 13326 22784 13670
rect 23768 13530 23796 16390
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 20916 11762 20944 12174
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21192 11558 21220 11698
rect 21468 11626 21496 12174
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21560 11558 21588 11766
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21192 11354 21220 11494
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21836 11286 21864 12174
rect 21928 11898 21956 12378
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 22756 11830 22784 13262
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 23860 9586 23888 16510
rect 24320 16454 24348 23054
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24780 22506 24808 22646
rect 24768 22500 24820 22506
rect 24768 22442 24820 22448
rect 25872 22500 25924 22506
rect 25872 22442 25924 22448
rect 25884 22098 25912 22442
rect 26068 22234 26096 27338
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26160 25702 26188 26318
rect 26252 26246 26280 27814
rect 26712 27470 26740 29650
rect 27264 29578 27292 30670
rect 27252 29572 27304 29578
rect 27252 29514 27304 29520
rect 27356 29510 27384 31146
rect 27540 30122 27568 31690
rect 27620 30728 27672 30734
rect 27620 30670 27672 30676
rect 27528 30116 27580 30122
rect 27528 30058 27580 30064
rect 27632 30054 27660 30670
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27344 29504 27396 29510
rect 27344 29446 27396 29452
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 26344 26314 26372 26726
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 26252 25974 26280 26182
rect 26344 26042 26372 26250
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26240 25968 26292 25974
rect 26240 25910 26292 25916
rect 26332 25832 26384 25838
rect 26332 25774 26384 25780
rect 26148 25696 26200 25702
rect 26148 25638 26200 25644
rect 26344 24954 26372 25774
rect 26332 24948 26384 24954
rect 26332 24890 26384 24896
rect 26344 24614 26372 24890
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26344 23186 26372 23462
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 25872 22092 25924 22098
rect 25872 22034 25924 22040
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24400 21956 24452 21962
rect 24400 21898 24452 21904
rect 24412 21690 24440 21898
rect 24872 21690 24900 21966
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24872 21146 24900 21626
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24492 19712 24544 19718
rect 24492 19654 24544 19660
rect 24504 19378 24532 19654
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24964 17610 24992 18702
rect 25792 18358 25820 19314
rect 25884 18358 25912 22034
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26252 21010 26280 21830
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26252 20466 26280 20946
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26344 19854 26372 20742
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 25976 18834 26004 19314
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25780 18352 25832 18358
rect 25780 18294 25832 18300
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 25976 18170 26004 18770
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 25884 18142 26004 18170
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 25332 16114 25360 17070
rect 25320 16108 25372 16114
rect 25320 16050 25372 16056
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24872 13326 24900 14282
rect 24964 14006 24992 14962
rect 25700 14074 25728 17546
rect 25884 16658 25912 18142
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 25976 17678 26004 18022
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 26068 17338 26096 18294
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 26056 17128 26108 17134
rect 26160 17082 26188 17546
rect 26252 17134 26280 19178
rect 26436 17678 26464 27270
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 26804 25838 26832 26522
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26516 25696 26568 25702
rect 26516 25638 26568 25644
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26528 25362 26556 25638
rect 26516 25356 26568 25362
rect 26516 25298 26568 25304
rect 26620 25294 26648 25638
rect 26608 25288 26660 25294
rect 26608 25230 26660 25236
rect 26792 25220 26844 25226
rect 26792 25162 26844 25168
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26528 24410 26556 24754
rect 26712 24410 26740 24822
rect 26804 24750 26832 25162
rect 26792 24744 26844 24750
rect 26792 24686 26844 24692
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26700 24404 26752 24410
rect 26700 24346 26752 24352
rect 26804 24274 26832 24686
rect 26884 24608 26936 24614
rect 26884 24550 26936 24556
rect 26792 24268 26844 24274
rect 26792 24210 26844 24216
rect 26804 23254 26832 24210
rect 26896 24206 26924 24550
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 26988 23730 27016 28018
rect 27356 27470 27384 29446
rect 27632 28626 27660 29990
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27724 28506 27752 30330
rect 27816 30258 27844 31826
rect 28276 31822 28304 32846
rect 29000 32836 29052 32842
rect 29000 32778 29052 32784
rect 28540 32496 28592 32502
rect 28540 32438 28592 32444
rect 28552 32026 28580 32438
rect 29012 32434 29040 32778
rect 30576 32502 30604 34682
rect 32324 33522 32352 34954
rect 32508 34474 32536 37198
rect 32680 37188 32732 37194
rect 32680 37130 32732 37136
rect 32692 35290 32720 37130
rect 33060 35630 33088 37266
rect 34164 35894 34192 39200
rect 34808 37346 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35346 37496 35402 37505
rect 35346 37431 35402 37440
rect 34808 37318 34928 37346
rect 35360 37330 35388 37431
rect 34900 36718 34928 37318
rect 35348 37324 35400 37330
rect 35348 37266 35400 37272
rect 34612 36712 34664 36718
rect 34612 36654 34664 36660
rect 34796 36712 34848 36718
rect 34796 36654 34848 36660
rect 34888 36712 34940 36718
rect 34888 36654 34940 36660
rect 34164 35866 34560 35894
rect 33048 35624 33100 35630
rect 33048 35566 33100 35572
rect 32680 35284 32732 35290
rect 32680 35226 32732 35232
rect 33692 35216 33744 35222
rect 33692 35158 33744 35164
rect 33600 35080 33652 35086
rect 33600 35022 33652 35028
rect 33612 34610 33640 35022
rect 33600 34604 33652 34610
rect 33600 34546 33652 34552
rect 32496 34468 32548 34474
rect 32496 34410 32548 34416
rect 32404 33924 32456 33930
rect 32404 33866 32456 33872
rect 32416 33658 32444 33866
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 30564 32496 30616 32502
rect 30564 32438 30616 32444
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 29092 32360 29144 32366
rect 29092 32302 29144 32308
rect 28724 32292 28776 32298
rect 28724 32234 28776 32240
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28736 31822 28764 32234
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28080 31748 28132 31754
rect 28080 31690 28132 31696
rect 28092 31482 28120 31690
rect 28080 31476 28132 31482
rect 28080 31418 28132 31424
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27896 29572 27948 29578
rect 27896 29514 27948 29520
rect 27632 28478 27752 28506
rect 27436 27532 27488 27538
rect 27436 27474 27488 27480
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27356 26382 27384 26930
rect 27448 26586 27476 27474
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27540 26926 27568 27406
rect 27632 26994 27660 28478
rect 27804 28416 27856 28422
rect 27804 28358 27856 28364
rect 27816 27606 27844 28358
rect 27804 27600 27856 27606
rect 27804 27542 27856 27548
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27528 26920 27580 26926
rect 27528 26862 27580 26868
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 27068 26240 27120 26246
rect 27068 26182 27120 26188
rect 27080 25294 27108 26182
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 27252 25288 27304 25294
rect 27252 25230 27304 25236
rect 27264 24886 27292 25230
rect 27252 24880 27304 24886
rect 27252 24822 27304 24828
rect 27356 24818 27384 26318
rect 27540 26042 27568 26862
rect 27620 26512 27672 26518
rect 27620 26454 27672 26460
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27632 25974 27660 26454
rect 27620 25968 27672 25974
rect 27620 25910 27672 25916
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27632 24750 27660 25774
rect 27724 25498 27752 27406
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27816 25906 27844 26522
rect 27908 26382 27936 29514
rect 28184 28762 28212 31214
rect 28276 30938 28304 31758
rect 28908 31272 28960 31278
rect 28908 31214 28960 31220
rect 28920 30938 28948 31214
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28908 30932 28960 30938
rect 28908 30874 28960 30880
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28644 30258 28672 30602
rect 28632 30252 28684 30258
rect 28632 30194 28684 30200
rect 28644 29850 28672 30194
rect 29000 30048 29052 30054
rect 29000 29990 29052 29996
rect 28632 29844 28684 29850
rect 28632 29786 28684 29792
rect 28172 28756 28224 28762
rect 28172 28698 28224 28704
rect 28184 28234 28212 28698
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28092 28206 28212 28234
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 28000 26586 28028 27542
rect 27988 26580 28040 26586
rect 27988 26522 28040 26528
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27804 25900 27856 25906
rect 27804 25842 27856 25848
rect 27712 25492 27764 25498
rect 27712 25434 27764 25440
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26792 23248 26844 23254
rect 26792 23190 26844 23196
rect 26988 23118 27016 23666
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 27356 22098 27384 24142
rect 27804 23792 27856 23798
rect 27804 23734 27856 23740
rect 27344 22092 27396 22098
rect 27816 22094 27844 23734
rect 27908 23526 27936 26318
rect 28000 24818 28028 26522
rect 28092 25838 28120 28206
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28080 25832 28132 25838
rect 28080 25774 28132 25780
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28000 24206 28028 24754
rect 28092 24342 28120 24754
rect 28184 24750 28212 28018
rect 28552 27606 28580 28494
rect 28540 27600 28592 27606
rect 28540 27542 28592 27548
rect 28644 26382 28672 29786
rect 29012 29578 29040 29990
rect 29000 29572 29052 29578
rect 29000 29514 29052 29520
rect 29012 28558 29040 29514
rect 29104 29510 29132 32302
rect 31116 32224 31168 32230
rect 31116 32166 31168 32172
rect 31128 32026 31156 32166
rect 31116 32020 31168 32026
rect 31116 31962 31168 31968
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 29748 30394 29776 31758
rect 30104 31748 30156 31754
rect 30104 31690 30156 31696
rect 30116 31482 30144 31690
rect 30104 31476 30156 31482
rect 30104 31418 30156 31424
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 29736 30388 29788 30394
rect 29736 30330 29788 30336
rect 29828 30252 29880 30258
rect 29828 30194 29880 30200
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 29840 29850 29868 30194
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 29828 29844 29880 29850
rect 29828 29786 29880 29792
rect 29932 29646 29960 29990
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29920 29640 29972 29646
rect 29920 29582 29972 29588
rect 29092 29504 29144 29510
rect 29092 29446 29144 29452
rect 29000 28552 29052 28558
rect 29000 28494 29052 28500
rect 29104 28218 29132 29446
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 29104 27470 29132 28154
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 29748 26994 29776 29582
rect 30024 29170 30052 30194
rect 30576 29850 30604 31282
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30668 29510 30696 30262
rect 31128 30258 31156 31962
rect 31116 30252 31168 30258
rect 31116 30194 31168 30200
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 30932 30048 30984 30054
rect 30932 29990 30984 29996
rect 30944 29714 30972 29990
rect 31128 29730 31156 30194
rect 30932 29708 30984 29714
rect 30932 29650 30984 29656
rect 31036 29702 31156 29730
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 30024 28626 30052 29106
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 30392 28642 30420 29038
rect 30012 28620 30064 28626
rect 30012 28562 30064 28568
rect 30300 28614 30420 28642
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30208 28082 30236 28494
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30208 27470 30236 28018
rect 30196 27464 30248 27470
rect 30196 27406 30248 27412
rect 29736 26988 29788 26994
rect 29736 26930 29788 26936
rect 29276 26920 29328 26926
rect 29276 26862 29328 26868
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 28632 26376 28684 26382
rect 28632 26318 28684 26324
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 28276 25906 28304 26318
rect 28264 25900 28316 25906
rect 28264 25842 28316 25848
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 28632 24608 28684 24614
rect 28632 24550 28684 24556
rect 28080 24336 28132 24342
rect 28080 24278 28132 24284
rect 28644 24274 28672 24550
rect 28920 24410 28948 24754
rect 29012 24682 29040 26318
rect 29092 26240 29144 26246
rect 29092 26182 29144 26188
rect 29104 25974 29132 26182
rect 29092 25968 29144 25974
rect 29092 25910 29144 25916
rect 29092 25288 29144 25294
rect 29092 25230 29144 25236
rect 29104 24818 29132 25230
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29000 24676 29052 24682
rect 29000 24618 29052 24624
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 28632 24268 28684 24274
rect 28632 24210 28684 24216
rect 27988 24200 28040 24206
rect 27988 24142 28040 24148
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28000 23662 28028 24142
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 27896 23520 27948 23526
rect 27896 23462 27948 23468
rect 27816 22066 27936 22094
rect 27344 22034 27396 22040
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27172 21622 27200 21966
rect 27724 21690 27752 21966
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27160 21616 27212 21622
rect 27160 21558 27212 21564
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 26712 21010 26740 21490
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26608 20868 26660 20874
rect 26608 20810 26660 20816
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26528 20058 26556 20402
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26620 19922 26648 20810
rect 26712 20534 26740 20946
rect 26700 20528 26752 20534
rect 26700 20470 26752 20476
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26988 19854 27016 20198
rect 27172 19854 27200 21558
rect 27724 21554 27752 21626
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27448 18902 27476 21286
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27724 19990 27752 20878
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27436 18896 27488 18902
rect 27436 18838 27488 18844
rect 27448 18442 27476 18838
rect 27264 18414 27476 18442
rect 26516 18284 26568 18290
rect 26516 18226 26568 18232
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26344 17338 26372 17614
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 26108 17076 26188 17082
rect 26056 17070 26188 17076
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26068 17054 26188 17070
rect 26160 16998 26188 17054
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 25976 16658 26004 16934
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25884 15366 25912 16594
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 26528 14346 26556 18226
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27172 18086 27200 18158
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27172 17678 27200 18022
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27172 17202 27200 17478
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27264 15978 27292 18414
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27448 17882 27476 18226
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 27252 15972 27304 15978
rect 27252 15914 27304 15920
rect 26700 15564 26752 15570
rect 26700 15506 26752 15512
rect 26712 15094 26740 15506
rect 27264 15502 27292 15914
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27264 15144 27292 15438
rect 27172 15116 27292 15144
rect 27356 15144 27384 16934
rect 27448 16046 27476 17138
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27448 15570 27476 15982
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27356 15116 27476 15144
rect 26700 15088 26752 15094
rect 26700 15030 26752 15036
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 25136 13932 25188 13938
rect 25136 13874 25188 13880
rect 25148 13530 25176 13874
rect 25700 13530 25728 14010
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 25700 12850 25728 13466
rect 26344 13190 26372 14214
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26804 12986 26832 13262
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 27172 12782 27200 15116
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27264 14618 27292 14962
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 27448 14414 27476 15116
rect 27540 14634 27568 19790
rect 27632 19378 27660 19790
rect 27620 19372 27672 19378
rect 27620 19314 27672 19320
rect 27632 18766 27660 19314
rect 27816 19258 27844 21830
rect 27908 20874 27936 22066
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 28000 21146 28028 21490
rect 28276 21457 28304 24142
rect 29104 23798 29132 24754
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29196 23866 29224 24142
rect 29184 23860 29236 23866
rect 29184 23802 29236 23808
rect 29092 23792 29144 23798
rect 29092 23734 29144 23740
rect 29288 22574 29316 26862
rect 29748 26314 29776 26930
rect 30300 26586 30328 28614
rect 30380 28484 30432 28490
rect 30380 28426 30432 28432
rect 30392 28014 30420 28426
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30392 27538 30420 27950
rect 30380 27532 30432 27538
rect 30380 27474 30432 27480
rect 30668 27402 30696 29446
rect 30656 27396 30708 27402
rect 30656 27338 30708 27344
rect 30288 26580 30340 26586
rect 30288 26522 30340 26528
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 29748 24410 29776 24754
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 29736 24404 29788 24410
rect 29736 24346 29788 24352
rect 29748 23798 29776 24346
rect 30208 24206 30236 24686
rect 30196 24200 30248 24206
rect 30196 24142 30248 24148
rect 30300 24070 30328 26522
rect 30748 25900 30800 25906
rect 30748 25842 30800 25848
rect 30380 25492 30432 25498
rect 30380 25434 30432 25440
rect 30288 24064 30340 24070
rect 30288 24006 30340 24012
rect 29736 23792 29788 23798
rect 29736 23734 29788 23740
rect 30392 23186 30420 25434
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30564 24948 30616 24954
rect 30564 24890 30616 24896
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30392 22642 30420 23122
rect 30576 22778 30604 24890
rect 30668 24818 30696 25094
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30668 24274 30696 24754
rect 30656 24268 30708 24274
rect 30656 24210 30708 24216
rect 30656 23588 30708 23594
rect 30656 23530 30708 23536
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 28262 21448 28318 21457
rect 28262 21383 28318 21392
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27908 19990 27936 20334
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 28000 20058 28028 20198
rect 27988 20052 28040 20058
rect 27988 19994 28040 20000
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 27988 19304 28040 19310
rect 27816 19230 27936 19258
rect 27988 19246 28040 19252
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27816 17882 27844 18226
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27632 16794 27660 17070
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27632 16658 27660 16730
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27632 16114 27660 16594
rect 27908 16454 27936 19230
rect 28000 18290 28028 19246
rect 28092 18902 28120 20402
rect 28080 18896 28132 18902
rect 28080 18838 28132 18844
rect 28184 18426 28212 20810
rect 28276 18834 28304 21383
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28460 20942 28488 21286
rect 28644 20942 28672 22170
rect 29564 21554 29592 22578
rect 30392 22522 30420 22578
rect 30392 22494 30512 22522
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 29644 21956 29696 21962
rect 29644 21898 29696 21904
rect 29656 21690 29684 21898
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 30392 21554 30420 22374
rect 30484 22234 30512 22494
rect 30472 22228 30524 22234
rect 30472 22170 30524 22176
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 30380 21548 30432 21554
rect 30380 21490 30432 21496
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28264 18828 28316 18834
rect 28264 18770 28316 18776
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28172 18420 28224 18426
rect 28172 18362 28224 18368
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27896 16448 27948 16454
rect 27896 16390 27948 16396
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 28000 15638 28028 18226
rect 28276 17678 28304 18566
rect 28460 17678 28488 18702
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28552 17542 28580 18702
rect 28644 17814 28672 20878
rect 29564 19854 29592 21490
rect 30576 20602 30604 22714
rect 30668 22574 30696 23530
rect 30760 23118 30788 25842
rect 30944 23594 30972 29650
rect 31036 29646 31064 29702
rect 31024 29640 31076 29646
rect 31024 29582 31076 29588
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 31036 28082 31064 29106
rect 31024 28076 31076 28082
rect 31024 28018 31076 28024
rect 31036 27674 31064 28018
rect 31128 27878 31156 29702
rect 31588 29102 31616 30194
rect 32508 29578 32536 30194
rect 32312 29572 32364 29578
rect 32312 29514 32364 29520
rect 32496 29572 32548 29578
rect 32496 29514 32548 29520
rect 31576 29096 31628 29102
rect 31576 29038 31628 29044
rect 31392 28960 31444 28966
rect 31392 28902 31444 28908
rect 31404 28558 31432 28902
rect 31588 28694 31616 29038
rect 31576 28688 31628 28694
rect 31576 28630 31628 28636
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31116 27872 31168 27878
rect 31116 27814 31168 27820
rect 31024 27668 31076 27674
rect 31024 27610 31076 27616
rect 31128 27538 31156 27814
rect 31116 27532 31168 27538
rect 31116 27474 31168 27480
rect 31404 27470 31432 28494
rect 32324 28218 32352 29514
rect 32312 28212 32364 28218
rect 32312 28154 32364 28160
rect 31760 28076 31812 28082
rect 31760 28018 31812 28024
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31392 27464 31444 27470
rect 31392 27406 31444 27412
rect 31392 25696 31444 25702
rect 31392 25638 31444 25644
rect 31404 25294 31432 25638
rect 31496 25294 31524 27814
rect 31680 27674 31708 27950
rect 31772 27946 31800 28018
rect 31760 27940 31812 27946
rect 31760 27882 31812 27888
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31772 27402 31800 27882
rect 32508 27538 32536 29514
rect 32692 29306 32720 30194
rect 33612 29850 33640 34546
rect 33704 33402 33732 35158
rect 33784 34400 33836 34406
rect 33784 34342 33836 34348
rect 33796 33590 33824 34342
rect 33876 34060 33928 34066
rect 33876 34002 33928 34008
rect 33784 33584 33836 33590
rect 33784 33526 33836 33532
rect 33888 33454 33916 34002
rect 34532 33454 34560 35866
rect 34624 35290 34652 36654
rect 34704 35624 34756 35630
rect 34704 35566 34756 35572
rect 34612 35284 34664 35290
rect 34612 35226 34664 35232
rect 34716 34202 34744 35566
rect 34808 35290 34836 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35348 35760 35400 35766
rect 35348 35702 35400 35708
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 35284 34848 35290
rect 34796 35226 34848 35232
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34704 34196 34756 34202
rect 34704 34138 34756 34144
rect 35360 33658 35388 35702
rect 35452 34066 35480 39200
rect 36912 37256 36964 37262
rect 36912 37198 36964 37204
rect 35806 36816 35862 36825
rect 35806 36751 35862 36760
rect 35820 35894 35848 36751
rect 35728 35866 35848 35894
rect 35728 34542 35756 35866
rect 35808 35624 35860 35630
rect 35808 35566 35860 35572
rect 35820 35290 35848 35566
rect 36728 35488 36780 35494
rect 36728 35430 36780 35436
rect 35808 35284 35860 35290
rect 35808 35226 35860 35232
rect 36740 34678 36768 35430
rect 36728 34672 36780 34678
rect 36728 34614 36780 34620
rect 35716 34536 35768 34542
rect 35716 34478 35768 34484
rect 36924 34202 36952 37198
rect 37188 36576 37240 36582
rect 37188 36518 37240 36524
rect 37200 36242 37228 36518
rect 37384 36310 37412 39200
rect 37832 37664 37884 37670
rect 38028 37618 38056 39200
rect 38290 38856 38346 38865
rect 38290 38791 38346 38800
rect 37832 37606 37884 37612
rect 37464 36848 37516 36854
rect 37464 36790 37516 36796
rect 37372 36304 37424 36310
rect 37372 36246 37424 36252
rect 37188 36236 37240 36242
rect 37188 36178 37240 36184
rect 37280 35012 37332 35018
rect 37280 34954 37332 34960
rect 36912 34196 36964 34202
rect 36912 34138 36964 34144
rect 35440 34060 35492 34066
rect 35440 34002 35492 34008
rect 36452 33992 36504 33998
rect 36452 33934 36504 33940
rect 35348 33652 35400 33658
rect 35348 33594 35400 33600
rect 36464 33590 36492 33934
rect 36820 33924 36872 33930
rect 36820 33866 36872 33872
rect 36832 33658 36860 33866
rect 36820 33652 36872 33658
rect 36820 33594 36872 33600
rect 36452 33584 36504 33590
rect 36452 33526 36504 33532
rect 33876 33448 33928 33454
rect 33704 33374 33824 33402
rect 33876 33390 33928 33396
rect 34520 33448 34572 33454
rect 34520 33390 34572 33396
rect 33796 31822 33824 33374
rect 33784 31816 33836 31822
rect 33784 31758 33836 31764
rect 33600 29844 33652 29850
rect 33600 29786 33652 29792
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 32496 27532 32548 27538
rect 32496 27474 32548 27480
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 31772 27062 31800 27338
rect 31760 27056 31812 27062
rect 31760 26998 31812 27004
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 31852 25424 31904 25430
rect 31852 25366 31904 25372
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 31404 24818 31432 25230
rect 31496 24954 31524 25230
rect 31484 24948 31536 24954
rect 31484 24890 31536 24896
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 31128 24138 31156 24754
rect 31116 24132 31168 24138
rect 31116 24074 31168 24080
rect 30932 23588 30984 23594
rect 30932 23530 30984 23536
rect 31864 23118 31892 25366
rect 30748 23112 30800 23118
rect 30748 23054 30800 23060
rect 31852 23112 31904 23118
rect 31852 23054 31904 23060
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31036 22642 31064 22918
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 30656 22568 30708 22574
rect 30656 22510 30708 22516
rect 30668 22094 30696 22510
rect 30668 22066 30788 22094
rect 30564 20596 30616 20602
rect 30564 20538 30616 20544
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29932 19854 29960 20198
rect 30104 19916 30156 19922
rect 30104 19858 30156 19864
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 28632 17808 28684 17814
rect 28632 17750 28684 17756
rect 29000 17808 29052 17814
rect 29000 17750 29052 17756
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 28368 16658 28396 16934
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28276 15978 28304 16526
rect 28264 15972 28316 15978
rect 28264 15914 28316 15920
rect 27988 15632 28040 15638
rect 27988 15574 28040 15580
rect 28276 15366 28304 15914
rect 28724 15904 28776 15910
rect 28724 15846 28776 15852
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 27540 14618 27660 14634
rect 27540 14612 27672 14618
rect 27540 14606 27620 14612
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27448 12782 27476 14350
rect 27540 13530 27568 14606
rect 27620 14554 27672 14560
rect 27896 14408 27948 14414
rect 27896 14350 27948 14356
rect 27908 14074 27936 14350
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27632 12850 27660 13126
rect 27816 12986 27844 13262
rect 28000 13190 28028 13874
rect 28736 13870 28764 15846
rect 29012 14618 29040 17750
rect 29104 15570 29132 19790
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29840 19446 29868 19654
rect 30116 19514 30144 19858
rect 30104 19508 30156 19514
rect 30104 19450 30156 19456
rect 29828 19440 29880 19446
rect 29828 19382 29880 19388
rect 30484 19174 30512 20402
rect 30760 20262 30788 22066
rect 33612 21554 33640 26318
rect 33796 23202 33824 31758
rect 33888 31278 33916 33390
rect 36360 33380 36412 33386
rect 36360 33322 36412 33328
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 36372 32858 36400 33322
rect 36452 33312 36504 33318
rect 36452 33254 36504 33260
rect 36464 32978 36492 33254
rect 36452 32972 36504 32978
rect 36452 32914 36504 32920
rect 36372 32830 36492 32858
rect 36464 32434 36492 32830
rect 36636 32836 36688 32842
rect 36636 32778 36688 32784
rect 36648 32570 36676 32778
rect 36636 32564 36688 32570
rect 36636 32506 36688 32512
rect 36452 32428 36504 32434
rect 36452 32370 36504 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35714 32056 35770 32065
rect 35714 31991 35770 32000
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34072 31414 34100 31622
rect 35728 31414 35756 31991
rect 34060 31408 34112 31414
rect 34060 31350 34112 31356
rect 35716 31408 35768 31414
rect 35716 31350 35768 31356
rect 33876 31272 33928 31278
rect 33876 31214 33928 31220
rect 33888 26518 33916 31214
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35256 28552 35308 28558
rect 35256 28494 35308 28500
rect 35268 28218 35296 28494
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 36004 28218 36032 28426
rect 35256 28212 35308 28218
rect 35256 28154 35308 28160
rect 35992 28212 36044 28218
rect 35992 28154 36044 28160
rect 36464 28082 36492 32370
rect 37188 29708 37240 29714
rect 37188 29650 37240 29656
rect 37200 28665 37228 29650
rect 37186 28656 37242 28665
rect 37186 28591 37242 28600
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 36452 27872 36504 27878
rect 36452 27814 36504 27820
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 36464 27538 36492 27814
rect 36452 27532 36504 27538
rect 36452 27474 36504 27480
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33876 26512 33928 26518
rect 33876 26454 33928 26460
rect 33888 23730 33916 26454
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 37292 24818 37320 34954
rect 37476 34610 37504 36790
rect 37648 36168 37700 36174
rect 37648 36110 37700 36116
rect 37660 35154 37688 36110
rect 37844 35894 37872 37606
rect 37752 35866 37872 35894
rect 37936 37590 38056 37618
rect 37648 35148 37700 35154
rect 37648 35090 37700 35096
rect 37556 35012 37608 35018
rect 37556 34954 37608 34960
rect 37568 34746 37596 34954
rect 37556 34740 37608 34746
rect 37556 34682 37608 34688
rect 37660 34626 37688 35090
rect 37464 34604 37516 34610
rect 37464 34546 37516 34552
rect 37568 34598 37688 34626
rect 37476 33522 37504 34546
rect 37464 33516 37516 33522
rect 37464 33458 37516 33464
rect 37372 33448 37424 33454
rect 37372 33390 37424 33396
rect 37280 24812 37332 24818
rect 37280 24754 37332 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35714 23896 35770 23905
rect 35714 23831 35770 23840
rect 35728 23798 35756 23831
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 33876 23724 33928 23730
rect 33876 23666 33928 23672
rect 34060 23656 34112 23662
rect 34060 23598 34112 23604
rect 34072 23322 34100 23598
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34060 23316 34112 23322
rect 34060 23258 34112 23264
rect 35438 23216 35494 23225
rect 33796 23174 33916 23202
rect 33888 23118 33916 23174
rect 35438 23151 35494 23160
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 30840 20324 30892 20330
rect 30840 20266 30892 20272
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 30748 20256 30800 20262
rect 30748 20198 30800 20204
rect 30472 19168 30524 19174
rect 30472 19110 30524 19116
rect 30484 18850 30512 19110
rect 30392 18822 30512 18850
rect 30392 18358 30420 18822
rect 30472 18692 30524 18698
rect 30472 18634 30524 18640
rect 30380 18352 30432 18358
rect 30380 18294 30432 18300
rect 30484 18290 30512 18634
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 30484 17882 30512 18226
rect 30472 17876 30524 17882
rect 30472 17818 30524 17824
rect 30288 17536 30340 17542
rect 30288 17478 30340 17484
rect 30300 17338 30328 17478
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30104 17196 30156 17202
rect 30104 17138 30156 17144
rect 30116 16454 30144 17138
rect 30300 16538 30328 17274
rect 30380 17196 30432 17202
rect 30380 17138 30432 17144
rect 30392 16794 30420 17138
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30472 16720 30524 16726
rect 30472 16662 30524 16668
rect 30484 16572 30512 16662
rect 30208 16510 30328 16538
rect 30392 16544 30512 16572
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30116 16114 30144 16390
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30012 16040 30064 16046
rect 30208 15994 30236 16510
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30300 16182 30328 16390
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 30392 16046 30420 16544
rect 30380 16040 30432 16046
rect 30064 15988 30328 15994
rect 30012 15982 30328 15988
rect 30380 15982 30432 15988
rect 30024 15966 30328 15982
rect 30196 15904 30248 15910
rect 30196 15846 30248 15852
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 29104 14958 29132 15506
rect 30104 15360 30156 15366
rect 30104 15302 30156 15308
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 29828 14340 29880 14346
rect 29828 14282 29880 14288
rect 29840 13938 29868 14282
rect 30116 14278 30144 15302
rect 30208 14958 30236 15846
rect 30300 15026 30328 15966
rect 30392 15502 30420 15982
rect 30576 15638 30604 20198
rect 30852 20074 30880 20266
rect 30760 20046 30880 20074
rect 30656 19780 30708 19786
rect 30656 19722 30708 19728
rect 30668 19378 30696 19722
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 30668 18902 30696 19314
rect 30656 18896 30708 18902
rect 30656 18838 30708 18844
rect 30760 17678 30788 20046
rect 30944 19394 30972 20538
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31128 20058 31156 20402
rect 31668 20392 31720 20398
rect 31668 20334 31720 20340
rect 31576 20324 31628 20330
rect 31576 20266 31628 20272
rect 31116 20052 31168 20058
rect 31116 19994 31168 20000
rect 31588 19854 31616 20266
rect 31680 20058 31708 20334
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31852 19916 31904 19922
rect 31852 19858 31904 19864
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 30852 19366 30972 19394
rect 30748 17672 30800 17678
rect 30748 17614 30800 17620
rect 30564 15632 30616 15638
rect 30564 15574 30616 15580
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30668 15162 30696 15438
rect 30852 15366 30880 19366
rect 30932 19304 30984 19310
rect 30932 19246 30984 19252
rect 30944 18290 30972 19246
rect 31864 18970 31892 19858
rect 31852 18964 31904 18970
rect 31852 18906 31904 18912
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 31680 18426 31708 18702
rect 31668 18420 31720 18426
rect 31668 18362 31720 18368
rect 32508 18290 32536 18702
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 31484 18284 31536 18290
rect 31484 18226 31536 18232
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 30944 17626 30972 18226
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 31208 18080 31260 18086
rect 31208 18022 31260 18028
rect 31128 17746 31156 18022
rect 31220 17814 31248 18022
rect 31208 17808 31260 17814
rect 31208 17750 31260 17756
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 31496 17678 31524 18226
rect 32048 17882 32076 18226
rect 32036 17876 32088 17882
rect 32036 17818 32088 17824
rect 31484 17672 31536 17678
rect 30944 17610 31064 17626
rect 31484 17614 31536 17620
rect 30944 17604 31076 17610
rect 30944 17598 31024 17604
rect 30944 16590 30972 17598
rect 31024 17546 31076 17552
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 30944 15978 30972 16526
rect 31312 16114 31340 16526
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 30932 15972 30984 15978
rect 30932 15914 30984 15920
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30288 15020 30340 15026
rect 30288 14962 30340 14968
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30104 14272 30156 14278
rect 30104 14214 30156 14220
rect 30116 13938 30144 14214
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28092 13326 28120 13806
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27160 12776 27212 12782
rect 27160 12718 27212 12724
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 27816 12238 27844 12922
rect 28000 12442 28028 13126
rect 29196 12918 29224 13874
rect 29920 13864 29972 13870
rect 29920 13806 29972 13812
rect 29932 13258 29960 13806
rect 29920 13252 29972 13258
rect 29920 13194 29972 13200
rect 29184 12912 29236 12918
rect 29184 12854 29236 12860
rect 28080 12640 28132 12646
rect 28080 12582 28132 12588
rect 27988 12436 28040 12442
rect 27988 12378 28040 12384
rect 28092 12238 28120 12582
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 29092 9444 29144 9450
rect 29092 9386 29144 9392
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19444 3998 19564 4026
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17224 2304 17276 2310
rect 17420 2258 17448 2314
rect 17512 2310 17540 2450
rect 17276 2252 17448 2258
rect 17224 2246 17448 2252
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17236 2230 17448 2246
rect 19352 800 19380 3334
rect 19444 3058 19472 3878
rect 19536 3398 19564 3998
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3602 20760 3878
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3126 20024 3470
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2926
rect 20824 2446 20852 5646
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 2650 20944 3402
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21284 800 21312 3538
rect 22020 3058 22048 3878
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24320 3058 24348 3470
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 22020 2446 22048 2858
rect 22204 2650 22232 2926
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22572 800 22600 2926
rect 23204 2916 23256 2922
rect 23204 2858 23256 2864
rect 23216 800 23244 2858
rect 24412 1850 24440 3334
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 2650 24532 2926
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 24596 2514 24624 3470
rect 24872 2514 24900 3878
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24964 2310 24992 4082
rect 25884 3602 25912 4558
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 26068 3602 26096 3878
rect 29104 3602 29132 9386
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 26056 3596 26108 3602
rect 26056 3538 26108 3544
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 24412 1822 24532 1850
rect 24504 800 24532 1822
rect 25148 800 25176 2450
rect 26436 800 26464 3538
rect 28264 3528 28316 3534
rect 28264 3470 28316 3476
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3126 28120 3334
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 27896 2984 27948 2990
rect 27896 2926 27948 2932
rect 27908 2650 27936 2926
rect 27896 2644 27948 2650
rect 27896 2586 27948 2592
rect 28276 2378 28304 3470
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 28368 800 28396 2926
rect 29932 2514 29960 13194
rect 32968 10062 32996 21490
rect 33888 17066 33916 23054
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 21622 35480 23151
rect 37186 22536 37242 22545
rect 37186 22471 37242 22480
rect 37200 22098 37228 22471
rect 37188 22092 37240 22098
rect 37188 22034 37240 22040
rect 35440 21616 35492 21622
rect 35440 21558 35492 21564
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 36452 18080 36504 18086
rect 36452 18022 36504 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 36464 17746 36492 18022
rect 36452 17740 36504 17746
rect 36452 17682 36504 17688
rect 37292 17202 37320 24754
rect 37384 19854 37412 33390
rect 37568 32314 37596 34598
rect 37648 34536 37700 34542
rect 37648 34478 37700 34484
rect 37660 32434 37688 34478
rect 37648 32428 37700 32434
rect 37648 32370 37700 32376
rect 37568 32286 37688 32314
rect 37660 30258 37688 32286
rect 37648 30252 37700 30258
rect 37648 30194 37700 30200
rect 37660 29238 37688 30194
rect 37648 29232 37700 29238
rect 37648 29174 37700 29180
rect 37556 27396 37608 27402
rect 37556 27338 37608 27344
rect 37568 27130 37596 27338
rect 37556 27124 37608 27130
rect 37556 27066 37608 27072
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37372 19848 37424 19854
rect 37372 19790 37424 19796
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 33876 17060 33928 17066
rect 33876 17002 33928 17008
rect 32956 10056 33008 10062
rect 32956 9998 33008 10004
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 30024 3602 30052 3878
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 33888 3534 33916 17002
rect 36636 16992 36688 16998
rect 36636 16934 36688 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 36648 16658 36676 16934
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36636 15904 36688 15910
rect 36636 15846 36688 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 36648 15570 36676 15846
rect 36636 15564 36688 15570
rect 36636 15506 36688 15512
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 37186 13016 37242 13025
rect 37186 12951 37242 12960
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 37200 12306 37228 12951
rect 37188 12300 37240 12306
rect 37188 12242 37240 12248
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 37188 11212 37240 11218
rect 37188 11154 37240 11160
rect 37200 10985 37228 11154
rect 37186 10976 37242 10985
rect 37186 10911 37242 10920
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34532 8945 34560 9454
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8968 34848 8974
rect 34518 8936 34574 8945
rect 34796 8910 34848 8916
rect 34518 8871 34574 8880
rect 34808 3942 34836 8910
rect 37186 8256 37242 8265
rect 34934 8188 35242 8197
rect 37186 8191 37242 8200
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 37200 7954 37228 8191
rect 37188 7948 37240 7954
rect 37188 7890 37240 7896
rect 37186 7576 37242 7585
rect 37186 7511 37242 7520
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 37200 6866 37228 7511
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37292 6322 37320 17138
rect 37384 16454 37412 19790
rect 37372 16448 37424 16454
rect 37372 16390 37424 16396
rect 37384 11762 37412 16390
rect 37476 15706 37504 22578
rect 37556 17604 37608 17610
rect 37556 17546 37608 17552
rect 37568 17338 37596 17546
rect 37556 17332 37608 17338
rect 37556 17274 37608 17280
rect 37660 16574 37688 29174
rect 37752 28626 37780 35866
rect 37936 35562 37964 37590
rect 38304 37330 38332 38791
rect 38292 37324 38344 37330
rect 38292 37266 38344 37272
rect 38016 37256 38068 37262
rect 38016 37198 38068 37204
rect 37924 35556 37976 35562
rect 37924 35498 37976 35504
rect 37832 35148 37884 35154
rect 37832 35090 37884 35096
rect 37844 34785 37872 35090
rect 37830 34776 37886 34785
rect 37830 34711 37886 34720
rect 37924 34672 37976 34678
rect 37924 34614 37976 34620
rect 37832 30796 37884 30802
rect 37832 30738 37884 30744
rect 37844 30705 37872 30738
rect 37830 30696 37886 30705
rect 37830 30631 37886 30640
rect 37740 28620 37792 28626
rect 37740 28562 37792 28568
rect 37936 28558 37964 34614
rect 37924 28552 37976 28558
rect 37924 28494 37976 28500
rect 37740 28484 37792 28490
rect 37740 28426 37792 28432
rect 37752 22642 37780 28426
rect 37832 25356 37884 25362
rect 37832 25298 37884 25304
rect 37844 25265 37872 25298
rect 37830 25256 37886 25265
rect 37830 25191 37886 25200
rect 37830 24576 37886 24585
rect 37830 24511 37886 24520
rect 37844 24274 37872 24511
rect 37832 24268 37884 24274
rect 37832 24210 37884 24216
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 37830 19136 37886 19145
rect 37830 19071 37886 19080
rect 37844 18834 37872 19071
rect 37832 18828 37884 18834
rect 37832 18770 37884 18776
rect 37660 16546 37780 16574
rect 37752 16114 37780 16546
rect 37740 16108 37792 16114
rect 37740 16050 37792 16056
rect 37648 15904 37700 15910
rect 37648 15846 37700 15852
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 37660 15638 37688 15846
rect 37648 15632 37700 15638
rect 37648 15574 37700 15580
rect 37372 11756 37424 11762
rect 37372 11698 37424 11704
rect 37556 7812 37608 7818
rect 37556 7754 37608 7760
rect 37568 7546 37596 7754
rect 37556 7540 37608 7546
rect 37556 7482 37608 7488
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37280 6316 37332 6322
rect 37280 6258 37332 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36912 5024 36964 5030
rect 36912 4966 36964 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35808 4072 35860 4078
rect 35808 4014 35860 4020
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 33980 3058 34008 3878
rect 34808 3534 34836 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 34060 3460 34112 3466
rect 34060 3402 34112 3408
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 29920 2508 29972 2514
rect 29920 2450 29972 2456
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 29012 800 29040 2382
rect 30932 2372 30984 2378
rect 30932 2314 30984 2320
rect 30944 800 30972 2314
rect 34072 1850 34100 3402
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 34164 3126 34192 3334
rect 34152 3120 34204 3126
rect 34152 3062 34204 3068
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34072 1822 34192 1850
rect 34164 800 34192 1822
rect 34808 800 34836 2926
rect 35820 2825 35848 4014
rect 36268 3596 36320 3602
rect 36268 3538 36320 3544
rect 36280 3058 36308 3538
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 35806 2816 35862 2825
rect 34934 2748 35242 2757
rect 35806 2751 35862 2760
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36924 2514 36952 4966
rect 37096 4684 37148 4690
rect 37096 4626 37148 4632
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 37108 2145 37136 4626
rect 37384 3670 37412 7346
rect 37752 6914 37780 16050
rect 37936 12850 37964 28494
rect 38028 23769 38056 37198
rect 38200 37188 38252 37194
rect 38200 37130 38252 37136
rect 38212 36922 38240 37130
rect 38672 37126 38700 39200
rect 39316 37670 39344 39200
rect 39304 37664 39356 37670
rect 39304 37606 39356 37612
rect 38660 37120 38712 37126
rect 38660 37062 38712 37068
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 38200 35692 38252 35698
rect 38200 35634 38252 35640
rect 38212 35222 38240 35634
rect 38200 35216 38252 35222
rect 38200 35158 38252 35164
rect 38108 30660 38160 30666
rect 38108 30602 38160 30608
rect 38120 30394 38148 30602
rect 38108 30388 38160 30394
rect 38108 30330 38160 30336
rect 38108 29572 38160 29578
rect 38108 29514 38160 29520
rect 38120 28762 38148 29514
rect 38108 28756 38160 28762
rect 38108 28698 38160 28704
rect 38212 28490 38240 35158
rect 38292 35080 38344 35086
rect 38292 35022 38344 35028
rect 38304 34610 38332 35022
rect 38292 34604 38344 34610
rect 38292 34546 38344 34552
rect 38290 34096 38346 34105
rect 38290 34031 38292 34040
rect 38344 34031 38346 34040
rect 38292 34002 38344 34008
rect 38290 33416 38346 33425
rect 38290 33351 38346 33360
rect 38304 32978 38332 33351
rect 38292 32972 38344 32978
rect 38292 32914 38344 32920
rect 38292 31136 38344 31142
rect 38292 31078 38344 31084
rect 38304 30802 38332 31078
rect 38292 30796 38344 30802
rect 38292 30738 38344 30744
rect 38384 29844 38436 29850
rect 38384 29786 38436 29792
rect 38292 29640 38344 29646
rect 38292 29582 38344 29588
rect 38304 29170 38332 29582
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38200 28484 38252 28490
rect 38200 28426 38252 28432
rect 38292 27396 38344 27402
rect 38292 27338 38344 27344
rect 38304 27305 38332 27338
rect 38290 27296 38346 27305
rect 38290 27231 38346 27240
rect 38396 25906 38424 29786
rect 38384 25900 38436 25906
rect 38384 25842 38436 25848
rect 38108 25696 38160 25702
rect 38108 25638 38160 25644
rect 38292 25696 38344 25702
rect 38292 25638 38344 25644
rect 38120 25362 38148 25638
rect 38304 25362 38332 25638
rect 38108 25356 38160 25362
rect 38108 25298 38160 25304
rect 38292 25356 38344 25362
rect 38292 25298 38344 25304
rect 38108 24608 38160 24614
rect 38108 24550 38160 24556
rect 38292 24608 38344 24614
rect 38292 24550 38344 24556
rect 38120 24274 38148 24550
rect 38304 24274 38332 24550
rect 38108 24268 38160 24274
rect 38108 24210 38160 24216
rect 38292 24268 38344 24274
rect 38292 24210 38344 24216
rect 38014 23760 38070 23769
rect 38014 23695 38070 23704
rect 38292 23112 38344 23118
rect 38292 23054 38344 23060
rect 38108 22432 38160 22438
rect 38108 22374 38160 22380
rect 38120 22098 38148 22374
rect 38304 22098 38332 23054
rect 38108 22092 38160 22098
rect 38108 22034 38160 22040
rect 38292 22092 38344 22098
rect 38292 22034 38344 22040
rect 38108 19712 38160 19718
rect 38108 19654 38160 19660
rect 38120 18834 38148 19654
rect 38292 19168 38344 19174
rect 38292 19110 38344 19116
rect 38304 18834 38332 19110
rect 38108 18828 38160 18834
rect 38108 18770 38160 18776
rect 38292 18828 38344 18834
rect 38292 18770 38344 18776
rect 38290 17776 38346 17785
rect 38290 17711 38292 17720
rect 38344 17711 38346 17720
rect 38292 17682 38344 17688
rect 38016 17196 38068 17202
rect 38016 17138 38068 17144
rect 38028 16794 38056 17138
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 38016 16788 38068 16794
rect 38016 16730 38068 16736
rect 37924 12844 37976 12850
rect 37924 12786 37976 12792
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37844 7954 37872 8230
rect 37832 7948 37884 7954
rect 37832 7890 37884 7896
rect 38028 7410 38056 16730
rect 38120 16726 38148 16934
rect 38108 16720 38160 16726
rect 38108 16662 38160 16668
rect 38304 16658 38332 17031
rect 38292 16652 38344 16658
rect 38292 16594 38344 16600
rect 38290 16416 38346 16425
rect 38290 16351 38346 16360
rect 38304 15570 38332 16351
rect 38292 15564 38344 15570
rect 38292 15506 38344 15512
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38108 12640 38160 12646
rect 38108 12582 38160 12588
rect 38120 12306 38148 12582
rect 38304 12306 38332 13262
rect 38108 12300 38160 12306
rect 38108 12242 38160 12248
rect 38292 12300 38344 12306
rect 38292 12242 38344 12248
rect 38108 11552 38160 11558
rect 38108 11494 38160 11500
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38120 11218 38148 11494
rect 38304 11218 38332 11494
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 38292 11212 38344 11218
rect 38292 11154 38344 11160
rect 38292 8968 38344 8974
rect 38292 8910 38344 8916
rect 38016 7404 38068 7410
rect 38016 7346 38068 7352
rect 38108 7200 38160 7206
rect 38108 7142 38160 7148
rect 37660 6886 37780 6914
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37476 3942 37504 4082
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37372 3664 37424 3670
rect 37372 3606 37424 3612
rect 37476 3058 37504 3878
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37188 2576 37240 2582
rect 37188 2518 37240 2524
rect 37094 2136 37150 2145
rect 37094 2071 37150 2080
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 5786 200 5898 800
rect 6430 200 6542 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10294 200 10406 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12226 200 12338 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 18666 200 18778 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21242 200 21354 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25106 200 25218 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 31546 200 31658 800
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 33478 200 33590 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
rect 36054 200 36166 800
rect 37200 105 37228 2518
rect 37660 2514 37688 6886
rect 38120 6866 38148 7142
rect 38304 6866 38332 8910
rect 38108 6860 38160 6866
rect 38108 6802 38160 6808
rect 38292 6860 38344 6866
rect 38292 6802 38344 6808
rect 38108 6112 38160 6118
rect 38108 6054 38160 6060
rect 38120 5778 38148 6054
rect 39304 5840 39356 5846
rect 39304 5782 39356 5788
rect 38108 5772 38160 5778
rect 38108 5714 38160 5720
rect 38292 5704 38344 5710
rect 38292 5646 38344 5652
rect 38304 5234 38332 5646
rect 38292 5228 38344 5234
rect 38292 5170 38344 5176
rect 38200 4616 38252 4622
rect 38200 4558 38252 4564
rect 38016 4548 38068 4554
rect 38016 4490 38068 4496
rect 38028 3194 38056 4490
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 38212 3058 38240 4558
rect 38660 3460 38712 3466
rect 38660 3402 38712 3408
rect 38200 3052 38252 3058
rect 38200 2994 38252 3000
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 38672 800 38700 3402
rect 39316 800 39344 5782
rect 37342 200 37454 800
rect 37986 200 38098 800
rect 38630 200 38742 800
rect 39274 200 39386 800
rect 37186 96 37242 105
rect 37186 31 37242 40
<< via2 >>
rect 1858 37440 1914 37496
rect 2778 38120 2834 38176
rect 1582 29280 1638 29336
rect 1858 22516 1860 22536
rect 1860 22516 1912 22536
rect 1912 22516 1914 22536
rect 1858 22480 1914 22516
rect 1582 21120 1638 21176
rect 1950 20476 1952 20496
rect 1952 20476 2004 20496
rect 2004 20476 2006 20496
rect 1950 20440 2006 20476
rect 1858 17076 1860 17096
rect 1860 17076 1912 17096
rect 1912 17076 1914 17096
rect 1858 17040 1914 17076
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 2778 33396 2780 33416
rect 2780 33396 2832 33416
rect 2832 33396 2834 33416
rect 2778 33360 2834 33396
rect 2778 30640 2834 30696
rect 3054 29960 3110 30016
rect 2870 28600 2926 28656
rect 2778 27956 2780 27976
rect 2780 27956 2832 27976
rect 2832 27956 2834 27976
rect 2778 27920 2834 27956
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 2778 21800 2834 21856
rect 2778 17720 2834 17776
rect 1582 8900 1638 8936
rect 1582 8880 1584 8900
rect 1584 8880 1636 8900
rect 1636 8880 1638 8900
rect 1582 8200 1638 8256
rect 1582 6860 1638 6896
rect 1582 6840 1584 6860
rect 1584 6840 1636 6860
rect 1636 6840 1638 6860
rect 1674 3440 1730 3496
rect 2778 15000 2834 15056
rect 2870 14320 2926 14376
rect 2778 12300 2834 12336
rect 2778 12280 2780 12300
rect 2780 12280 2832 12300
rect 2832 12280 2834 12300
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 26560 4122 26616
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1858 2372 1914 2408
rect 1858 2352 1860 2372
rect 1860 2352 1912 2372
rect 1912 2352 1914 2372
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4066 19796 4068 19816
rect 4068 19796 4120 19816
rect 4120 19796 4122 19816
rect 4066 19760 4122 19796
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12960 4122 13016
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3054 2760 3110 2816
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2962 2080 3018 2136
rect 2870 1400 2926 1456
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 10598 22616 10654 22672
rect 10690 18844 10692 18864
rect 10692 18844 10744 18864
rect 10744 18844 10746 18864
rect 10690 18808 10746 18844
rect 14462 19660 14464 19680
rect 14464 19660 14516 19680
rect 14516 19660 14518 19680
rect 14462 19624 14518 19660
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 12622 11348 12678 11384
rect 12622 11328 12624 11348
rect 12624 11328 12676 11348
rect 12676 11328 12678 11348
rect 17222 20884 17224 20904
rect 17224 20884 17276 20904
rect 17276 20884 17278 20904
rect 17222 20848 17278 20884
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19890 33360 19946 33416
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20442 33360 20498 33416
rect 21178 33360 21234 33416
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 17866 18808 17922 18864
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20718 22636 20774 22672
rect 20718 22616 20720 22636
rect 20720 22616 20772 22636
rect 20772 22616 20774 22636
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 18878 19624 18934 19680
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 20902 23740 20904 23760
rect 20904 23740 20956 23760
rect 20956 23740 20958 23760
rect 20902 23704 20958 23740
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 18510 11328 18566 11384
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 21914 21412 21970 21448
rect 21914 21392 21916 21412
rect 21916 21392 21968 21412
rect 21968 21392 21970 21412
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35346 37440 35402 37496
rect 28262 21392 28318 21448
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35806 36760 35862 36816
rect 38290 38800 38346 38856
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35714 32000 35770 32056
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 37186 28600 37242 28656
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35714 23840 35770 23896
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35438 23160 35494 23216
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 37186 22480 37242 22536
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 37186 12960 37242 13016
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37186 10920 37242 10976
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34518 8880 34574 8936
rect 37186 8200 37242 8256
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 37186 7520 37242 7576
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37830 34720 37886 34776
rect 37830 30640 37886 30696
rect 37830 25200 37886 25256
rect 37830 24520 37886 24576
rect 37830 19080 37886 19136
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35806 2760 35862 2816
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 34060 38346 34096
rect 38290 34040 38292 34060
rect 38292 34040 38344 34060
rect 38344 34040 38346 34060
rect 38290 33360 38346 33416
rect 38290 27240 38346 27296
rect 38014 23704 38070 23760
rect 38290 17740 38346 17776
rect 38290 17720 38292 17740
rect 38292 17720 38344 17740
rect 38344 17720 38346 17740
rect 38290 17040 38346 17096
rect 38290 16360 38346 16416
rect 37094 2080 37150 2136
rect 2778 720 2834 776
rect 37186 40 37242 96
<< metal3 >>
rect 200 39388 800 39628
rect 39200 39388 39800 39628
rect 38285 38858 38351 38861
rect 39200 38858 39800 38948
rect 38285 38856 39800 38858
rect 38285 38800 38290 38856
rect 38346 38800 39800 38856
rect 38285 38798 39800 38800
rect 38285 38795 38351 38798
rect 39200 38708 39800 38798
rect 200 38178 800 38268
rect 2773 38178 2839 38181
rect 200 38176 2839 38178
rect 200 38120 2778 38176
rect 2834 38120 2839 38176
rect 200 38118 2839 38120
rect 200 38028 800 38118
rect 2773 38115 2839 38118
rect 39200 38028 39800 38268
rect 200 37498 800 37588
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 1853 37498 1919 37501
rect 200 37496 1919 37498
rect 200 37440 1858 37496
rect 1914 37440 1919 37496
rect 200 37438 1919 37440
rect 200 37348 800 37438
rect 1853 37435 1919 37438
rect 35341 37498 35407 37501
rect 39200 37498 39800 37588
rect 35341 37496 39800 37498
rect 35341 37440 35346 37496
rect 35402 37440 39800 37496
rect 35341 37438 39800 37440
rect 35341 37435 35407 37438
rect 39200 37348 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36668 800 36908
rect 35801 36818 35867 36821
rect 39200 36818 39800 36908
rect 35801 36816 39800 36818
rect 35801 36760 35806 36816
rect 35862 36760 39800 36816
rect 35801 36758 39800 36760
rect 35801 36755 35867 36758
rect 39200 36668 39800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 35988 800 36228
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35308 800 35548
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 39200 35308 39800 35548
rect 200 34628 800 34868
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 37825 34778 37891 34781
rect 39200 34778 39800 34868
rect 37825 34776 39800 34778
rect 37825 34720 37830 34776
rect 37886 34720 39800 34776
rect 37825 34718 39800 34720
rect 37825 34715 37891 34718
rect 39200 34628 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 33948 800 34188
rect 38285 34098 38351 34101
rect 39200 34098 39800 34188
rect 38285 34096 39800 34098
rect 38285 34040 38290 34096
rect 38346 34040 39800 34096
rect 38285 34038 39800 34040
rect 38285 34035 38351 34038
rect 39200 33948 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33508
rect 2773 33418 2839 33421
rect 200 33416 2839 33418
rect 200 33360 2778 33416
rect 2834 33360 2839 33416
rect 200 33358 2839 33360
rect 200 33268 800 33358
rect 2773 33355 2839 33358
rect 19885 33418 19951 33421
rect 20437 33418 20503 33421
rect 21173 33418 21239 33421
rect 19885 33416 21239 33418
rect 19885 33360 19890 33416
rect 19946 33360 20442 33416
rect 20498 33360 21178 33416
rect 21234 33360 21239 33416
rect 19885 33358 21239 33360
rect 19885 33355 19951 33358
rect 20437 33355 20503 33358
rect 21173 33355 21239 33358
rect 38285 33418 38351 33421
rect 39200 33418 39800 33508
rect 38285 33416 39800 33418
rect 38285 33360 38290 33416
rect 38346 33360 39800 33416
rect 38285 33358 39800 33360
rect 38285 33355 38351 33358
rect 39200 33268 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32588 800 32828
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 39200 32588 39800 32828
rect 200 31908 800 32148
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 35709 32058 35775 32061
rect 39200 32058 39800 32148
rect 35709 32056 39800 32058
rect 35709 32000 35714 32056
rect 35770 32000 39800 32056
rect 35709 31998 39800 32000
rect 35709 31995 35775 31998
rect 39200 31908 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 39200 31228 39800 31468
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30788
rect 2773 30698 2839 30701
rect 200 30696 2839 30698
rect 200 30640 2778 30696
rect 2834 30640 2839 30696
rect 200 30638 2839 30640
rect 200 30548 800 30638
rect 2773 30635 2839 30638
rect 37825 30698 37891 30701
rect 39200 30698 39800 30788
rect 37825 30696 39800 30698
rect 37825 30640 37830 30696
rect 37886 30640 39800 30696
rect 37825 30638 39800 30640
rect 37825 30635 37891 30638
rect 39200 30548 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 200 30018 800 30108
rect 3049 30018 3115 30021
rect 200 30016 3115 30018
rect 200 29960 3054 30016
rect 3110 29960 3115 30016
rect 200 29958 3115 29960
rect 200 29868 800 29958
rect 3049 29955 3115 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 39200 29868 39800 30108
rect 200 29338 800 29428
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1577 29338 1643 29341
rect 200 29336 1643 29338
rect 200 29280 1582 29336
rect 1638 29280 1643 29336
rect 200 29278 1643 29280
rect 200 29188 800 29278
rect 1577 29275 1643 29278
rect 39200 29188 39800 29428
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28748
rect 2865 28658 2931 28661
rect 200 28656 2931 28658
rect 200 28600 2870 28656
rect 2926 28600 2931 28656
rect 200 28598 2931 28600
rect 200 28508 800 28598
rect 2865 28595 2931 28598
rect 37181 28658 37247 28661
rect 39200 28658 39800 28748
rect 37181 28656 39800 28658
rect 37181 28600 37186 28656
rect 37242 28600 39800 28656
rect 37181 28598 39800 28600
rect 37181 28595 37247 28598
rect 39200 28508 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 200 27978 800 28068
rect 2773 27978 2839 27981
rect 200 27976 2839 27978
rect 200 27920 2778 27976
rect 2834 27920 2839 27976
rect 200 27918 2839 27920
rect 200 27828 800 27918
rect 2773 27915 2839 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27148 800 27388
rect 38285 27298 38351 27301
rect 39200 27298 39800 27388
rect 38285 27296 39800 27298
rect 38285 27240 38290 27296
rect 38346 27240 39800 27296
rect 38285 27238 39800 27240
rect 38285 27235 38351 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 39200 27148 39800 27238
rect 200 26618 800 26708
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4061 26618 4127 26621
rect 200 26616 4127 26618
rect 200 26560 4066 26616
rect 4122 26560 4127 26616
rect 200 26558 4127 26560
rect 200 26468 800 26558
rect 4061 26555 4127 26558
rect 39200 26468 39800 26708
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25788 800 26028
rect 39200 25788 39800 26028
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25108 800 25348
rect 37825 25258 37891 25261
rect 39200 25258 39800 25348
rect 37825 25256 39800 25258
rect 37825 25200 37830 25256
rect 37886 25200 39800 25256
rect 37825 25198 39800 25200
rect 37825 25195 37891 25198
rect 39200 25108 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24428 800 24668
rect 37825 24578 37891 24581
rect 39200 24578 39800 24668
rect 37825 24576 39800 24578
rect 37825 24520 37830 24576
rect 37886 24520 39800 24576
rect 37825 24518 39800 24520
rect 37825 24515 37891 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 39200 24428 39800 24518
rect 200 23748 800 23988
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 35709 23898 35775 23901
rect 39200 23898 39800 23988
rect 35709 23896 39800 23898
rect 35709 23840 35714 23896
rect 35770 23840 39800 23896
rect 35709 23838 39800 23840
rect 35709 23835 35775 23838
rect 20897 23762 20963 23765
rect 38009 23762 38075 23765
rect 20897 23760 38075 23762
rect 20897 23704 20902 23760
rect 20958 23704 38014 23760
rect 38070 23704 38075 23760
rect 39200 23748 39800 23838
rect 20897 23702 38075 23704
rect 20897 23699 20963 23702
rect 38009 23699 38075 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 35433 23218 35499 23221
rect 39200 23218 39800 23308
rect 35433 23216 39800 23218
rect 35433 23160 35438 23216
rect 35494 23160 39800 23216
rect 35433 23158 39800 23160
rect 35433 23155 35499 23158
rect 39200 23068 39800 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 10593 22674 10659 22677
rect 20713 22674 20779 22677
rect 10593 22672 20779 22674
rect 200 22538 800 22628
rect 10593 22616 10598 22672
rect 10654 22616 20718 22672
rect 20774 22616 20779 22672
rect 10593 22614 20779 22616
rect 10593 22611 10659 22614
rect 20713 22611 20779 22614
rect 1853 22538 1919 22541
rect 200 22536 1919 22538
rect 200 22480 1858 22536
rect 1914 22480 1919 22536
rect 200 22478 1919 22480
rect 200 22388 800 22478
rect 1853 22475 1919 22478
rect 37181 22538 37247 22541
rect 39200 22538 39800 22628
rect 37181 22536 39800 22538
rect 37181 22480 37186 22536
rect 37242 22480 39800 22536
rect 37181 22478 39800 22480
rect 37181 22475 37247 22478
rect 39200 22388 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 200 21858 800 21948
rect 2773 21858 2839 21861
rect 200 21856 2839 21858
rect 200 21800 2778 21856
rect 2834 21800 2839 21856
rect 200 21798 2839 21800
rect 200 21708 800 21798
rect 2773 21795 2839 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 39200 21708 39800 21948
rect 21909 21450 21975 21453
rect 28257 21450 28323 21453
rect 21909 21448 28323 21450
rect 21909 21392 21914 21448
rect 21970 21392 28262 21448
rect 28318 21392 28323 21448
rect 21909 21390 28323 21392
rect 21909 21387 21975 21390
rect 28257 21387 28323 21390
rect 200 21178 800 21268
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1577 21178 1643 21181
rect 200 21176 1643 21178
rect 200 21120 1582 21176
rect 1638 21120 1643 21176
rect 200 21118 1643 21120
rect 200 21028 800 21118
rect 1577 21115 1643 21118
rect 39200 21028 39800 21268
rect 17217 20906 17283 20909
rect 17350 20906 17356 20908
rect 17217 20904 17356 20906
rect 17217 20848 17222 20904
rect 17278 20848 17356 20904
rect 17217 20846 17356 20848
rect 17217 20843 17283 20846
rect 17350 20844 17356 20846
rect 17420 20844 17426 20908
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20588
rect 1945 20498 2011 20501
rect 200 20496 2011 20498
rect 200 20440 1950 20496
rect 2006 20440 2011 20496
rect 200 20438 2011 20440
rect 200 20348 800 20438
rect 1945 20435 2011 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19908
rect 4061 19818 4127 19821
rect 200 19816 4127 19818
rect 200 19760 4066 19816
rect 4122 19760 4127 19816
rect 200 19758 4127 19760
rect 200 19668 800 19758
rect 4061 19755 4127 19758
rect 14457 19682 14523 19685
rect 18873 19682 18939 19685
rect 14457 19680 18939 19682
rect 14457 19624 14462 19680
rect 14518 19624 18878 19680
rect 18934 19624 18939 19680
rect 39200 19668 39800 19908
rect 14457 19622 18939 19624
rect 14457 19619 14523 19622
rect 18873 19619 18939 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 200 18988 800 19228
rect 37825 19138 37891 19141
rect 39200 19138 39800 19228
rect 37825 19136 39800 19138
rect 37825 19080 37830 19136
rect 37886 19080 39800 19136
rect 37825 19078 39800 19080
rect 37825 19075 37891 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 39200 18988 39800 19078
rect 10685 18866 10751 18869
rect 17861 18866 17927 18869
rect 10685 18864 17927 18866
rect 10685 18808 10690 18864
rect 10746 18808 17866 18864
rect 17922 18808 17927 18864
rect 10685 18806 17927 18808
rect 10685 18803 10751 18806
rect 17861 18803 17927 18806
rect 200 18308 800 18548
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 39200 18308 39800 18548
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17868
rect 2773 17778 2839 17781
rect 200 17776 2839 17778
rect 200 17720 2778 17776
rect 2834 17720 2839 17776
rect 200 17718 2839 17720
rect 200 17628 800 17718
rect 2773 17715 2839 17718
rect 38285 17778 38351 17781
rect 39200 17778 39800 17868
rect 38285 17776 39800 17778
rect 38285 17720 38290 17776
rect 38346 17720 39800 17776
rect 38285 17718 39800 17720
rect 38285 17715 38351 17718
rect 39200 17628 39800 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 200 17098 800 17188
rect 1853 17098 1919 17101
rect 200 17096 1919 17098
rect 200 17040 1858 17096
rect 1914 17040 1919 17096
rect 200 17038 1919 17040
rect 200 16948 800 17038
rect 1853 17035 1919 17038
rect 38285 17098 38351 17101
rect 39200 17098 39800 17188
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 16948 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 200 16268 800 16508
rect 38285 16418 38351 16421
rect 39200 16418 39800 16508
rect 38285 16416 39800 16418
rect 38285 16360 38290 16416
rect 38346 16360 39800 16416
rect 38285 16358 39800 16360
rect 38285 16355 38351 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 39200 16268 39800 16358
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 39200 15588 39800 15828
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 200 15058 800 15148
rect 2773 15058 2839 15061
rect 200 15056 2839 15058
rect 200 15000 2778 15056
rect 2834 15000 2839 15056
rect 200 14998 2839 15000
rect 200 14908 800 14998
rect 2773 14995 2839 14998
rect 39200 14908 39800 15148
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14468
rect 2865 14378 2931 14381
rect 200 14376 2931 14378
rect 200 14320 2870 14376
rect 2926 14320 2931 14376
rect 200 14318 2931 14320
rect 200 14228 800 14318
rect 2865 14315 2931 14318
rect 39200 14228 39800 14468
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13548 800 13788
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 39200 13548 39800 13788
rect 200 13018 800 13108
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4061 13018 4127 13021
rect 200 13016 4127 13018
rect 200 12960 4066 13016
rect 4122 12960 4127 13016
rect 200 12958 4127 12960
rect 200 12868 800 12958
rect 4061 12955 4127 12958
rect 37181 13018 37247 13021
rect 39200 13018 39800 13108
rect 37181 13016 39800 13018
rect 37181 12960 37186 13016
rect 37242 12960 39800 13016
rect 37181 12958 39800 12960
rect 37181 12955 37247 12958
rect 39200 12868 39800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12428
rect 2773 12338 2839 12341
rect 200 12336 2839 12338
rect 200 12280 2778 12336
rect 2834 12280 2839 12336
rect 200 12278 2839 12280
rect 200 12188 800 12278
rect 2773 12275 2839 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 200 11508 800 11748
rect 39200 11508 39800 11748
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 12617 11386 12683 11389
rect 18505 11386 18571 11389
rect 12617 11384 18571 11386
rect 12617 11328 12622 11384
rect 12678 11328 18510 11384
rect 18566 11328 18571 11384
rect 12617 11326 18571 11328
rect 12617 11323 12683 11326
rect 18505 11323 18571 11326
rect 200 10828 800 11068
rect 37181 10978 37247 10981
rect 39200 10978 39800 11068
rect 37181 10976 39800 10978
rect 37181 10920 37186 10976
rect 37242 10920 39800 10976
rect 37181 10918 39800 10920
rect 37181 10915 37247 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 39200 10828 39800 10918
rect 200 10148 800 10388
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 39200 10148 39800 10388
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9468 800 9708
rect 39200 9468 39800 9708
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 9028
rect 1577 8938 1643 8941
rect 200 8936 1643 8938
rect 200 8880 1582 8936
rect 1638 8880 1643 8936
rect 200 8878 1643 8880
rect 200 8788 800 8878
rect 1577 8875 1643 8878
rect 34513 8938 34579 8941
rect 39200 8938 39800 9028
rect 34513 8936 39800 8938
rect 34513 8880 34518 8936
rect 34574 8880 39800 8936
rect 34513 8878 39800 8880
rect 34513 8875 34579 8878
rect 39200 8788 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 200 8258 800 8348
rect 1577 8258 1643 8261
rect 200 8256 1643 8258
rect 200 8200 1582 8256
rect 1638 8200 1643 8256
rect 200 8198 1643 8200
rect 200 8108 800 8198
rect 1577 8195 1643 8198
rect 37181 8258 37247 8261
rect 39200 8258 39800 8348
rect 37181 8256 39800 8258
rect 37181 8200 37186 8256
rect 37242 8200 39800 8256
rect 37181 8198 39800 8200
rect 37181 8195 37247 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 39200 8108 39800 8198
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 37181 7578 37247 7581
rect 39200 7578 39800 7668
rect 37181 7576 39800 7578
rect 37181 7520 37186 7576
rect 37242 7520 39800 7576
rect 37181 7518 39800 7520
rect 37181 7515 37247 7518
rect 39200 7428 39800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6988
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6748 800 6838
rect 1577 6835 1643 6838
rect 39200 6748 39800 6988
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 200 6068 800 6308
rect 39200 6068 39800 6308
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5388 800 5628
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 39200 5388 39800 5628
rect 200 4708 800 4948
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 200 4028 800 4268
rect 39200 4028 39800 4268
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3588
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3348 800 3438
rect 1669 3435 1735 3438
rect 39200 3348 39800 3588
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2908
rect 3049 2818 3115 2821
rect 200 2816 3115 2818
rect 200 2760 3054 2816
rect 3110 2760 3115 2816
rect 200 2758 3115 2760
rect 200 2668 800 2758
rect 3049 2755 3115 2758
rect 35801 2818 35867 2821
rect 39200 2818 39800 2908
rect 35801 2816 39800 2818
rect 35801 2760 35806 2816
rect 35862 2760 39800 2816
rect 35801 2758 39800 2760
rect 35801 2755 35867 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 39200 2668 39800 2758
rect 1853 2410 1919 2413
rect 17350 2410 17356 2412
rect 1853 2408 17356 2410
rect 1853 2352 1858 2408
rect 1914 2352 17356 2408
rect 1853 2350 17356 2352
rect 1853 2347 1919 2350
rect 17350 2348 17356 2350
rect 17420 2348 17426 2412
rect 200 2138 800 2228
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 2957 2138 3023 2141
rect 200 2136 3023 2138
rect 200 2080 2962 2136
rect 3018 2080 3023 2136
rect 200 2078 3023 2080
rect 200 1988 800 2078
rect 2957 2075 3023 2078
rect 37089 2138 37155 2141
rect 39200 2138 39800 2228
rect 37089 2136 39800 2138
rect 37089 2080 37094 2136
rect 37150 2080 39800 2136
rect 37089 2078 39800 2080
rect 37089 2075 37155 2078
rect 39200 1988 39800 2078
rect 200 1458 800 1548
rect 2865 1458 2931 1461
rect 200 1456 2931 1458
rect 200 1400 2870 1456
rect 2926 1400 2931 1456
rect 200 1398 2931 1400
rect 200 1308 800 1398
rect 2865 1395 2931 1398
rect 39200 1308 39800 1548
rect 200 778 800 868
rect 2773 778 2839 781
rect 200 776 2839 778
rect 200 720 2778 776
rect 2834 720 2839 776
rect 200 718 2839 720
rect 200 628 800 718
rect 2773 715 2839 718
rect 39200 628 39800 868
rect 37181 98 37247 101
rect 39200 98 39800 188
rect 37181 96 39800 98
rect 37181 40 37186 96
rect 37242 40 39800 96
rect 37181 38 39800 40
rect 37181 35 37247 38
rect 39200 -52 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 17356 20844 17420 20908
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 17356 2348 17420 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 17355 20908 17421 20909
rect 17355 20844 17356 20908
rect 17420 20844 17421 20908
rect 17355 20843 17421 20844
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 17358 2413 17418 20843
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 17355 2412 17421 2413
rect 17355 2348 17356 2412
rect 17420 2348 17421 2412
rect 17355 2347 17421 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1667941163
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1667941163
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1667941163
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1667941163
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1667941163
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1667941163
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1667941163
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_236
timestamp 1667941163
transform 1 0 22816 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_240
timestamp 1667941163
transform 1 0 23184 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1667941163
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_289
timestamp 1667941163
transform 1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_295
timestamp 1667941163
transform 1 0 28244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1667941163
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1667941163
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1667941163
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1667941163
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1667941163
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_289
timestamp 1667941163
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_312
timestamp 1667941163
transform 1 0 29808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324
timestamp 1667941163
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_378
timestamp 1667941163
transform 1 0 35880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_398
timestamp 1667941163
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_36
timestamp 1667941163
transform 1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_43
timestamp 1667941163
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1667941163
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_69
timestamp 1667941163
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1667941163
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_122
timestamp 1667941163
transform 1 0 12328 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1667941163
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1667941163
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_204
timestamp 1667941163
transform 1 0 19872 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_212
timestamp 1667941163
transform 1 0 20608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_241
timestamp 1667941163
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1667941163
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_259
timestamp 1667941163
transform 1 0 24932 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_267
timestamp 1667941163
transform 1 0 25668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_290
timestamp 1667941163
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_297
timestamp 1667941163
transform 1 0 28428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1667941163
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1667941163
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_335
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_347
timestamp 1667941163
transform 1 0 33028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_355
timestamp 1667941163
transform 1 0 33764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1667941163
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_374
timestamp 1667941163
transform 1 0 35512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_399
timestamp 1667941163
transform 1 0 37812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1667941163
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_47
timestamp 1667941163
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1667941163
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_119
timestamp 1667941163
transform 1 0 12052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_131
timestamp 1667941163
transform 1 0 13156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_143
timestamp 1667941163
transform 1 0 14260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_155
timestamp 1667941163
transform 1 0 15364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_204
timestamp 1667941163
transform 1 0 19872 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_212
timestamp 1667941163
transform 1 0 20608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_230
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_242
timestamp 1667941163
transform 1 0 23368 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_254
timestamp 1667941163
transform 1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_260
timestamp 1667941163
transform 1 0 25024 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_268
timestamp 1667941163
transform 1 0 25760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_313
timestamp 1667941163
transform 1 0 29900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_360
timestamp 1667941163
transform 1 0 34224 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_368
timestamp 1667941163
transform 1 0 34960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1667941163
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_398
timestamp 1667941163
transform 1 0 37720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1667941163
transform 1 0 2392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1667941163
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_45
timestamp 1667941163
transform 1 0 5244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1667941163
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_69
timestamp 1667941163
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1667941163
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_269
timestamp 1667941163
transform 1 0 25852 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_273
timestamp 1667941163
transform 1 0 26220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_285
timestamp 1667941163
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1667941163
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_404
timestamp 1667941163
transform 1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1667941163
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1667941163
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1667941163
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1667941163
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1667941163
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_400
timestamp 1667941163
transform 1 0 37904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1667941163
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_12
timestamp 1667941163
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_19
timestamp 1667941163
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_383
timestamp 1667941163
transform 1 0 36340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1667941163
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_16
timestamp 1667941163
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_28
timestamp 1667941163
transform 1 0 3680 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_40
timestamp 1667941163
transform 1 0 4784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1667941163
transform 1 0 5336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1667941163
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_398
timestamp 1667941163
transform 1 0 37720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_406
timestamp 1667941163
transform 1 0 38456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1667941163
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_67
timestamp 1667941163
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1667941163
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_383
timestamp 1667941163
transform 1 0 36340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1667941163
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_12
timestamp 1667941163
transform 1 0 2208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1667941163
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_36
timestamp 1667941163
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_44
timestamp 1667941163
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1667941163
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_398
timestamp 1667941163
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_383
timestamp 1667941163
transform 1 0 36340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1667941163
transform 1 0 37904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1667941163
transform 1 0 38456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_400
timestamp 1667941163
transform 1 0 37904 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1667941163
transform 1 0 38456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1667941163
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1667941163
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_18
timestamp 1667941163
transform 1 0 2760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_30
timestamp 1667941163
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1667941163
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_243
timestamp 1667941163
transform 1 0 23460 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_268
timestamp 1667941163
transform 1 0 25760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_185
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1667941163
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1667941163
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_16
timestamp 1667941163
transform 1 0 2576 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1667941163
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1667941163
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_187
timestamp 1667941163
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_209
timestamp 1667941163
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1667941163
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1667941163
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1667941163
transform 1 0 11868 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1667941163
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_147
timestamp 1667941163
transform 1 0 14628 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_159
timestamp 1667941163
transform 1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_166
timestamp 1667941163
transform 1 0 16376 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_178
timestamp 1667941163
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1667941163
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_205
timestamp 1667941163
transform 1 0 19964 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_211
timestamp 1667941163
transform 1 0 20516 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_383
timestamp 1667941163
transform 1 0 36340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1667941163
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1667941163
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1667941163
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1667941163
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1667941163
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_99
timestamp 1667941163
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_120
timestamp 1667941163
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_132
timestamp 1667941163
transform 1 0 13248 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1667941163
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_157
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_177
timestamp 1667941163
transform 1 0 17388 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_201
timestamp 1667941163
transform 1 0 19596 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_209
timestamp 1667941163
transform 1 0 20332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_232
timestamp 1667941163
transform 1 0 22448 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_244
timestamp 1667941163
transform 1 0 23552 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_256
timestamp 1667941163
transform 1 0 24656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_268
timestamp 1667941163
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_398
timestamp 1667941163
transform 1 0 37720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1667941163
transform 1 0 10672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_112
timestamp 1667941163
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1667941163
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_130
timestamp 1667941163
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_152
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1667941163
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_178
timestamp 1667941163
transform 1 0 17480 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1667941163
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1667941163
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_211
timestamp 1667941163
transform 1 0 20516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1667941163
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_223
timestamp 1667941163
transform 1 0 21620 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_229
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_241
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1667941163
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_294
timestamp 1667941163
transform 1 0 28152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1667941163
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_383
timestamp 1667941163
transform 1 0 36340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_405
timestamp 1667941163
transform 1 0 38364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_13
timestamp 1667941163
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_25
timestamp 1667941163
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_37
timestamp 1667941163
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1667941163
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_92
timestamp 1667941163
transform 1 0 9568 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_98
timestamp 1667941163
transform 1 0 10120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_133
timestamp 1667941163
transform 1 0 13340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1667941163
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_158
timestamp 1667941163
transform 1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1667941163
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1667941163
transform 1 0 17848 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_190
timestamp 1667941163
transform 1 0 18584 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_196
timestamp 1667941163
transform 1 0 19136 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1667941163
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_210
timestamp 1667941163
transform 1 0 20424 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_249
timestamp 1667941163
transform 1 0 24012 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1667941163
transform 1 0 24748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_266
timestamp 1667941163
transform 1 0 25576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1667941163
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_291
timestamp 1667941163
transform 1 0 27876 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_301
timestamp 1667941163
transform 1 0 28796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_313
timestamp 1667941163
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1667941163
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_398
timestamp 1667941163
transform 1 0 37720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1667941163
transform 1 0 38456 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_117
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1667941163
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1667941163
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1667941163
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_184
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_225
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_231
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_238
timestamp 1667941163
transform 1 0 23000 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_244
timestamp 1667941163
transform 1 0 23552 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_262
timestamp 1667941163
transform 1 0 25208 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_270
timestamp 1667941163
transform 1 0 25944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_280
timestamp 1667941163
transform 1 0 26864 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_294
timestamp 1667941163
transform 1 0 28152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_400
timestamp 1667941163
transform 1 0 37904 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1667941163
transform 1 0 38456 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_14
timestamp 1667941163
transform 1 0 2392 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_26
timestamp 1667941163
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_38
timestamp 1667941163
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1667941163
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_100
timestamp 1667941163
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_121
timestamp 1667941163
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_128
timestamp 1667941163
transform 1 0 12880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1667941163
transform 1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_189
timestamp 1667941163
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_196
timestamp 1667941163
transform 1 0 19136 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_207
timestamp 1667941163
transform 1 0 20148 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_215
timestamp 1667941163
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_244
timestamp 1667941163
transform 1 0 23552 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_252
timestamp 1667941163
transform 1 0 24288 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1667941163
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_289
timestamp 1667941163
transform 1 0 27692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_298
timestamp 1667941163
transform 1 0 28520 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_302
timestamp 1667941163
transform 1 0 28888 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_308
timestamp 1667941163
transform 1 0 29440 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_322
timestamp 1667941163
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1667941163
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1667941163
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1667941163
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1667941163
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_116
timestamp 1667941163
transform 1 0 11776 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_128
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1667941163
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1667941163
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_218
timestamp 1667941163
transform 1 0 21160 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_226
timestamp 1667941163
transform 1 0 21896 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1667941163
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_283
timestamp 1667941163
transform 1 0 27140 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_292
timestamp 1667941163
transform 1 0 27968 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1667941163
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_316
timestamp 1667941163
transform 1 0 30176 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_328
timestamp 1667941163
transform 1 0 31280 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_340
timestamp 1667941163
transform 1 0 32384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_352
timestamp 1667941163
transform 1 0 33488 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_29
timestamp 1667941163
transform 1 0 3772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_41
timestamp 1667941163
transform 1 0 4876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1667941163
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1667941163
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_129
timestamp 1667941163
transform 1 0 12972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1667941163
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_140
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_144
timestamp 1667941163
transform 1 0 14352 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_156
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_200
timestamp 1667941163
transform 1 0 19504 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1667941163
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1667941163
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1667941163
transform 1 0 23460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_260
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1667941163
transform 1 0 25760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_313
timestamp 1667941163
transform 1 0 29900 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_322
timestamp 1667941163
transform 1 0 30728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1667941163
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_40
timestamp 1667941163
transform 1 0 4784 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_52
timestamp 1667941163
transform 1 0 5888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_64
timestamp 1667941163
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1667941163
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_89
timestamp 1667941163
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_166
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1667941163
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_184
timestamp 1667941163
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_203
timestamp 1667941163
transform 1 0 19780 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_227
timestamp 1667941163
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_241
timestamp 1667941163
transform 1 0 23276 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1667941163
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_261
timestamp 1667941163
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_279
timestamp 1667941163
transform 1 0 26772 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_290
timestamp 1667941163
transform 1 0 27784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_302
timestamp 1667941163
transform 1 0 28888 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1667941163
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_313
timestamp 1667941163
transform 1 0 29900 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_322
timestamp 1667941163
transform 1 0 30728 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_334
timestamp 1667941163
transform 1 0 31832 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_346
timestamp 1667941163
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1667941163
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_383
timestamp 1667941163
transform 1 0 36340 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_25
timestamp 1667941163
transform 1 0 3404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1667941163
transform 1 0 4784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1667941163
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_155
timestamp 1667941163
transform 1 0 15364 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1667941163
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1667941163
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_198
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_210
timestamp 1667941163
transform 1 0 20424 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_218
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_243
timestamp 1667941163
transform 1 0 23460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_255
timestamp 1667941163
transform 1 0 24564 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_268
timestamp 1667941163
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1667941163
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_307
timestamp 1667941163
transform 1 0 29348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_315
timestamp 1667941163
transform 1 0 30084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_322
timestamp 1667941163
transform 1 0 30728 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1667941163
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_400
timestamp 1667941163
transform 1 0 37904 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1667941163
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_12
timestamp 1667941163
transform 1 0 2208 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_37
timestamp 1667941163
transform 1 0 4508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_49
timestamp 1667941163
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_61
timestamp 1667941163
transform 1 0 6716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1667941163
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1667941163
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1667941163
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_98
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1667941163
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1667941163
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1667941163
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1667941163
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_149
timestamp 1667941163
transform 1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1667941163
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_163
timestamp 1667941163
transform 1 0 16100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_169
timestamp 1667941163
transform 1 0 16652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_173
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_182
timestamp 1667941163
transform 1 0 17848 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_229
timestamp 1667941163
transform 1 0 22172 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_241
timestamp 1667941163
transform 1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1667941163
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_278
timestamp 1667941163
transform 1 0 26680 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_290
timestamp 1667941163
transform 1 0 27784 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1667941163
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1667941163
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_322
timestamp 1667941163
transform 1 0 30728 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_329
timestamp 1667941163
transform 1 0 31372 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_341
timestamp 1667941163
transform 1 0 32476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_353
timestamp 1667941163
transform 1 0 33580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1667941163
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_383
timestamp 1667941163
transform 1 0 36340 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1667941163
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1667941163
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_41
timestamp 1667941163
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1667941163
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 1667941163
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_154
timestamp 1667941163
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1667941163
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1667941163
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_255
timestamp 1667941163
transform 1 0 24564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_264
timestamp 1667941163
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_288
timestamp 1667941163
transform 1 0 27600 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_300
timestamp 1667941163
transform 1 0 28704 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_312
timestamp 1667941163
transform 1 0 29808 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1667941163
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1667941163
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_398
timestamp 1667941163
transform 1 0 37720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_8
timestamp 1667941163
transform 1 0 1840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_22
timestamp 1667941163
transform 1 0 3128 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_37
timestamp 1667941163
transform 1 0 4508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_49
timestamp 1667941163
transform 1 0 5612 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_61
timestamp 1667941163
transform 1 0 6716 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_73
timestamp 1667941163
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1667941163
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_91
timestamp 1667941163
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_98
timestamp 1667941163
transform 1 0 10120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1667941163
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_114
timestamp 1667941163
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1667941163
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1667941163
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1667941163
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_178
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1667941163
transform 1 0 18032 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1667941163
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_276
timestamp 1667941163
transform 1 0 26496 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_284
timestamp 1667941163
transform 1 0 27232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_299
timestamp 1667941163
transform 1 0 28612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_317
timestamp 1667941163
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_327
timestamp 1667941163
transform 1 0 31188 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_337
timestamp 1667941163
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_349
timestamp 1667941163
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1667941163
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_383
timestamp 1667941163
transform 1 0 36340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_405
timestamp 1667941163
transform 1 0 38364 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1667941163
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_29
timestamp 1667941163
transform 1 0 3772 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1667941163
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_179
timestamp 1667941163
transform 1 0 17572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_187
timestamp 1667941163
transform 1 0 18308 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_194
timestamp 1667941163
transform 1 0 18952 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1667941163
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_234
timestamp 1667941163
transform 1 0 22632 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_246
timestamp 1667941163
transform 1 0 23736 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_258
timestamp 1667941163
transform 1 0 24840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1667941163
transform 1 0 25576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_288
timestamp 1667941163
transform 1 0 27600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_308
timestamp 1667941163
transform 1 0 29440 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_316
timestamp 1667941163
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_327
timestamp 1667941163
transform 1 0 31188 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1667941163
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_342
timestamp 1667941163
transform 1 0 32568 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_354
timestamp 1667941163
transform 1 0 33672 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_366
timestamp 1667941163
transform 1 0 34776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_378
timestamp 1667941163
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1667941163
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_398
timestamp 1667941163
transform 1 0 37720 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1667941163
transform 1 0 38456 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_13
timestamp 1667941163
transform 1 0 2300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1667941163
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_42
timestamp 1667941163
transform 1 0 4968 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_54
timestamp 1667941163
transform 1 0 6072 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_66
timestamp 1667941163
transform 1 0 7176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1667941163
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_92
timestamp 1667941163
transform 1 0 9568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_101
timestamp 1667941163
transform 1 0 10396 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_166
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_172
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_182
timestamp 1667941163
transform 1 0 17848 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1667941163
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_216
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1667941163
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_236
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1667941163
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_262
timestamp 1667941163
transform 1 0 25208 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_274
timestamp 1667941163
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1667941163
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_294
timestamp 1667941163
transform 1 0 28152 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1667941163
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_328
timestamp 1667941163
transform 1 0 31280 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_335
timestamp 1667941163
transform 1 0 31924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_347
timestamp 1667941163
transform 1 0 33028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1667941163
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_383
timestamp 1667941163
transform 1 0 36340 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_34
timestamp 1667941163
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1667941163
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_136
timestamp 1667941163
transform 1 0 13616 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_144
timestamp 1667941163
transform 1 0 14352 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_151
timestamp 1667941163
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1667941163
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_182
timestamp 1667941163
transform 1 0 17848 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_189
timestamp 1667941163
transform 1 0 18492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_201
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_207
timestamp 1667941163
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1667941163
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1667941163
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1667941163
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1667941163
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_255
timestamp 1667941163
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_267
timestamp 1667941163
transform 1 0 25668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_287
timestamp 1667941163
transform 1 0 27508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_299
timestamp 1667941163
transform 1 0 28612 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_330
timestamp 1667941163
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1667941163
transform 1 0 37904 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1667941163
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_12
timestamp 1667941163
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_19
timestamp 1667941163
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1667941163
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1667941163
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_166
timestamp 1667941163
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_170
timestamp 1667941163
transform 1 0 16744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1667941163
transform 1 0 17664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1667941163
transform 1 0 18216 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_205
timestamp 1667941163
transform 1 0 19964 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_222
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_234
timestamp 1667941163
transform 1 0 22632 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_242
timestamp 1667941163
transform 1 0 23368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_276
timestamp 1667941163
transform 1 0 26496 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_280
timestamp 1667941163
transform 1 0 26864 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1667941163
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_293
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1667941163
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_314
timestamp 1667941163
transform 1 0 29992 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_327
timestamp 1667941163
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_338
timestamp 1667941163
transform 1 0 32200 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_350
timestamp 1667941163
transform 1 0 33304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1667941163
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_398
timestamp 1667941163
transform 1 0 37720 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1667941163
transform 1 0 38456 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_30
timestamp 1667941163
transform 1 0 3864 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_42
timestamp 1667941163
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_88
timestamp 1667941163
transform 1 0 9200 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_95
timestamp 1667941163
transform 1 0 9844 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_121
timestamp 1667941163
transform 1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1667941163
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1667941163
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1667941163
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1667941163
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_235
timestamp 1667941163
transform 1 0 22724 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_247
timestamp 1667941163
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_259
timestamp 1667941163
transform 1 0 24932 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_267
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_288
timestamp 1667941163
transform 1 0 27600 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_296
timestamp 1667941163
transform 1 0 28336 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_308
timestamp 1667941163
transform 1 0 29440 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_316
timestamp 1667941163
transform 1 0 30176 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_326
timestamp 1667941163
transform 1 0 31096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1667941163
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_92
timestamp 1667941163
transform 1 0 9568 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_116
timestamp 1667941163
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_150
timestamp 1667941163
transform 1 0 14904 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_162
timestamp 1667941163
transform 1 0 16008 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_170
timestamp 1667941163
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_176
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1667941163
transform 1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1667941163
transform 1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_234
timestamp 1667941163
transform 1 0 22632 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1667941163
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1667941163
transform 1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1667941163
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_293
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_300
timestamp 1667941163
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_16
timestamp 1667941163
transform 1 0 2576 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_23
timestamp 1667941163
transform 1 0 3220 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_35
timestamp 1667941163
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1667941163
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1667941163
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_94
timestamp 1667941163
transform 1 0 9752 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_106
timestamp 1667941163
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_122
timestamp 1667941163
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1667941163
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_138
timestamp 1667941163
transform 1 0 13800 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1667941163
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_175
timestamp 1667941163
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_182
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_190
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_195
timestamp 1667941163
transform 1 0 19044 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_207
timestamp 1667941163
transform 1 0 20148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1667941163
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_239
timestamp 1667941163
transform 1 0 23092 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_245
timestamp 1667941163
transform 1 0 23644 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_254
timestamp 1667941163
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_312
timestamp 1667941163
transform 1 0 29808 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_324
timestamp 1667941163
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_345
timestamp 1667941163
transform 1 0 32844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_374
timestamp 1667941163
transform 1 0 35512 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1667941163
transform 1 0 36616 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_103
timestamp 1667941163
transform 1 0 10580 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1667941163
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_132
timestamp 1667941163
transform 1 0 13248 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_163
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_171
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_183
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_205
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_219
timestamp 1667941163
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_231
timestamp 1667941163
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_243
timestamp 1667941163
transform 1 0 23460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1667941163
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_257
timestamp 1667941163
transform 1 0 24748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_274
timestamp 1667941163
transform 1 0 26312 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1667941163
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1667941163
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_328
timestamp 1667941163
transform 1 0 31280 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_340
timestamp 1667941163
transform 1 0 32384 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_352
timestamp 1667941163
transform 1 0 33488 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_383
timestamp 1667941163
transform 1 0 36340 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 1667941163
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_29
timestamp 1667941163
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_41
timestamp 1667941163
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_90
timestamp 1667941163
transform 1 0 9384 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_102
timestamp 1667941163
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_121
timestamp 1667941163
transform 1 0 12236 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_128
timestamp 1667941163
transform 1 0 12880 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_140
timestamp 1667941163
transform 1 0 13984 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_157
timestamp 1667941163
transform 1 0 15548 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_176
timestamp 1667941163
transform 1 0 17296 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1667941163
transform 1 0 18032 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_194
timestamp 1667941163
transform 1 0 18952 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1667941163
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1667941163
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1667941163
transform 1 0 23644 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_253
timestamp 1667941163
transform 1 0 24380 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_260
timestamp 1667941163
transform 1 0 25024 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1667941163
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_326
timestamp 1667941163
transform 1 0 31096 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1667941163
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_398
timestamp 1667941163
transform 1 0 37720 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1667941163
transform 1 0 38456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_14
timestamp 1667941163
transform 1 0 2392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1667941163
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1667941163
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1667941163
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_104
timestamp 1667941163
transform 1 0 10672 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_122
timestamp 1667941163
transform 1 0 12328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_129
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1667941163
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_146
timestamp 1667941163
transform 1 0 14536 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1667941163
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_162
timestamp 1667941163
transform 1 0 16008 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_167
timestamp 1667941163
transform 1 0 16468 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_176
timestamp 1667941163
transform 1 0 17296 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_180
timestamp 1667941163
transform 1 0 17664 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_205
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_212
timestamp 1667941163
transform 1 0 20608 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_231
timestamp 1667941163
transform 1 0 22356 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_242
timestamp 1667941163
transform 1 0 23368 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1667941163
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_280
timestamp 1667941163
transform 1 0 26864 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_292
timestamp 1667941163
transform 1 0 27968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1667941163
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_317
timestamp 1667941163
transform 1 0 30268 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_326
timestamp 1667941163
transform 1 0 31096 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_337
timestamp 1667941163
transform 1 0 32108 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_349
timestamp 1667941163
transform 1 0 33212 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1667941163
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_400
timestamp 1667941163
transform 1 0 37904 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1667941163
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1667941163
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_100
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_124
timestamp 1667941163
transform 1 0 12512 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_179
timestamp 1667941163
transform 1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_203
timestamp 1667941163
transform 1 0 19780 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_209
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1667941163
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_231
timestamp 1667941163
transform 1 0 22356 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_239
timestamp 1667941163
transform 1 0 23092 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_247
timestamp 1667941163
transform 1 0 23828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_253
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_270
timestamp 1667941163
transform 1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1667941163
transform 1 0 28796 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_310
timestamp 1667941163
transform 1 0 29624 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_322
timestamp 1667941163
transform 1 0 30728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1667941163
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_355
timestamp 1667941163
transform 1 0 33764 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_377
timestamp 1667941163
transform 1 0 35788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1667941163
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_46
timestamp 1667941163
transform 1 0 5336 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_58
timestamp 1667941163
transform 1 0 6440 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_70
timestamp 1667941163
transform 1 0 7544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_78
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_93
timestamp 1667941163
transform 1 0 9660 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_99
timestamp 1667941163
transform 1 0 10212 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_116
timestamp 1667941163
transform 1 0 11776 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_124
timestamp 1667941163
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1667941163
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1667941163
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1667941163
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_164
timestamp 1667941163
transform 1 0 16192 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_168
timestamp 1667941163
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1667941163
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_205
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1667941163
transform 1 0 22080 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1667941163
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1667941163
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_262
timestamp 1667941163
transform 1 0 25208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_274
timestamp 1667941163
transform 1 0 26312 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_281
timestamp 1667941163
transform 1 0 26956 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1667941163
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_303
timestamp 1667941163
transform 1 0 28980 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_317
timestamp 1667941163
transform 1 0 30268 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_329
timestamp 1667941163
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_341
timestamp 1667941163
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1667941163
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1667941163
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_383
timestamp 1667941163
transform 1 0 36340 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1667941163
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_95
timestamp 1667941163
transform 1 0 9844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 1667941163
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_141
timestamp 1667941163
transform 1 0 14076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_182
timestamp 1667941163
transform 1 0 17848 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_189
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_201
timestamp 1667941163
transform 1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_207
timestamp 1667941163
transform 1 0 20148 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_214
timestamp 1667941163
transform 1 0 20792 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_255
timestamp 1667941163
transform 1 0 24564 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1667941163
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_289
timestamp 1667941163
transform 1 0 27692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_296
timestamp 1667941163
transform 1 0 28336 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1667941163
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_311
timestamp 1667941163
transform 1 0 29716 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_320
timestamp 1667941163
transform 1 0 30544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1667941163
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_398
timestamp 1667941163
transform 1 0 37720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_34
timestamp 1667941163
transform 1 0 4232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1667941163
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_58
timestamp 1667941163
transform 1 0 6440 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_70
timestamp 1667941163
transform 1 0 7544 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1667941163
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_125
timestamp 1667941163
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1667941163
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1667941163
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_155
timestamp 1667941163
transform 1 0 15364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_167
timestamp 1667941163
transform 1 0 16468 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1667941163
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1667941163
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_205
timestamp 1667941163
transform 1 0 19964 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_217
timestamp 1667941163
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_222
timestamp 1667941163
transform 1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_230
timestamp 1667941163
transform 1 0 22264 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1667941163
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_259
timestamp 1667941163
transform 1 0 24932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_271
timestamp 1667941163
transform 1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_279
timestamp 1667941163
transform 1 0 26772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_288
timestamp 1667941163
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_300
timestamp 1667941163
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_317
timestamp 1667941163
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_324
timestamp 1667941163
transform 1 0 30912 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_331
timestamp 1667941163
transform 1 0 31556 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_343
timestamp 1667941163
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_355
timestamp 1667941163
transform 1 0 33764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_383
timestamp 1667941163
transform 1 0 36340 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_86
timestamp 1667941163
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1667941163
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_122
timestamp 1667941163
transform 1 0 12328 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_139
timestamp 1667941163
transform 1 0 13892 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_147
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_155
timestamp 1667941163
transform 1 0 15364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1667941163
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1667941163
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_188
timestamp 1667941163
transform 1 0 18400 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1667941163
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_241
timestamp 1667941163
transform 1 0 23276 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_262
timestamp 1667941163
transform 1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_270
timestamp 1667941163
transform 1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_274
timestamp 1667941163
transform 1 0 26312 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1667941163
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_291
timestamp 1667941163
transform 1 0 27876 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_299
timestamp 1667941163
transform 1 0 28612 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_316
timestamp 1667941163
transform 1 0 30176 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1667941163
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_398
timestamp 1667941163
transform 1 0 37720 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_52
timestamp 1667941163
transform 1 0 5888 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_64
timestamp 1667941163
transform 1 0 6992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_76
timestamp 1667941163
transform 1 0 8096 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_94
timestamp 1667941163
transform 1 0 9752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_102
timestamp 1667941163
transform 1 0 10488 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_130
timestamp 1667941163
transform 1 0 13064 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_164
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_176
timestamp 1667941163
transform 1 0 17296 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_183
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_203
timestamp 1667941163
transform 1 0 19780 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_215
timestamp 1667941163
transform 1 0 20884 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_234
timestamp 1667941163
transform 1 0 22632 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_259
timestamp 1667941163
transform 1 0 24932 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_267
timestamp 1667941163
transform 1 0 25668 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_273
timestamp 1667941163
transform 1 0 26220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_282
timestamp 1667941163
transform 1 0 27048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_295
timestamp 1667941163
transform 1 0 28244 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_315
timestamp 1667941163
transform 1 0 30084 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_327
timestamp 1667941163
transform 1 0 31188 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_339
timestamp 1667941163
transform 1 0 32292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_351
timestamp 1667941163
transform 1 0 33396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_31
timestamp 1667941163
transform 1 0 3956 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_35
timestamp 1667941163
transform 1 0 4324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_47
timestamp 1667941163
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1667941163
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_91
timestamp 1667941163
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_103
timestamp 1667941163
transform 1 0 10580 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_122
timestamp 1667941163
transform 1 0 12328 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_128
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_140
timestamp 1667941163
transform 1 0 13984 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_152
timestamp 1667941163
transform 1 0 15088 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1667941163
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1667941163
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_187
timestamp 1667941163
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_199
timestamp 1667941163
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_211
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_248
timestamp 1667941163
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_255
timestamp 1667941163
transform 1 0 24564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_263
timestamp 1667941163
transform 1 0 25300 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_269
timestamp 1667941163
transform 1 0 25852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1667941163
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_319
timestamp 1667941163
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1667941163
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_398
timestamp 1667941163
transform 1 0 37720 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1667941163
transform 1 0 38456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_13
timestamp 1667941163
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1667941163
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_96
timestamp 1667941163
transform 1 0 9936 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_102
timestamp 1667941163
transform 1 0 10488 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_110
timestamp 1667941163
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_122
timestamp 1667941163
transform 1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_126
timestamp 1667941163
transform 1 0 12696 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1667941163
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_162
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_170
timestamp 1667941163
transform 1 0 16744 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_206
timestamp 1667941163
transform 1 0 20056 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_219
timestamp 1667941163
transform 1 0 21252 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_231
timestamp 1667941163
transform 1 0 22356 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_235
timestamp 1667941163
transform 1 0 22724 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_240
timestamp 1667941163
transform 1 0 23184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_264
timestamp 1667941163
transform 1 0 25392 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_276
timestamp 1667941163
transform 1 0 26496 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_282
timestamp 1667941163
transform 1 0 27048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_290
timestamp 1667941163
transform 1 0 27784 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1667941163
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 1667941163
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_323
timestamp 1667941163
transform 1 0 30820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_334
timestamp 1667941163
transform 1 0 31832 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_341
timestamp 1667941163
transform 1 0 32476 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1667941163
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1667941163
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_383
timestamp 1667941163
transform 1 0 36340 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_7
timestamp 1667941163
transform 1 0 1748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_29
timestamp 1667941163
transform 1 0 3772 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_38
timestamp 1667941163
transform 1 0 4600 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_50
timestamp 1667941163
transform 1 0 5704 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_89
timestamp 1667941163
transform 1 0 9292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_101
timestamp 1667941163
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1667941163
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_122
timestamp 1667941163
transform 1 0 12328 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_135
timestamp 1667941163
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_147
timestamp 1667941163
transform 1 0 14628 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_154
timestamp 1667941163
transform 1 0 15272 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_176
timestamp 1667941163
transform 1 0 17296 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_188
timestamp 1667941163
transform 1 0 18400 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1667941163
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_233
timestamp 1667941163
transform 1 0 22540 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_238
timestamp 1667941163
transform 1 0 23000 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1667941163
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_256
timestamp 1667941163
transform 1 0 24656 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1667941163
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_289
timestamp 1667941163
transform 1 0 27692 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_307
timestamp 1667941163
transform 1 0 29348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_319
timestamp 1667941163
transform 1 0 30452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1667941163
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_344
timestamp 1667941163
transform 1 0 32752 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_356
timestamp 1667941163
transform 1 0 33856 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_368
timestamp 1667941163
transform 1 0 34960 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_372
timestamp 1667941163
transform 1 0 35328 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1667941163
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1667941163
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_399
timestamp 1667941163
transform 1 0 37812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_12
timestamp 1667941163
transform 1 0 2208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_16
timestamp 1667941163
transform 1 0 2576 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1667941163
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 1667941163
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_55
timestamp 1667941163
transform 1 0 6164 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_67
timestamp 1667941163
transform 1 0 7268 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_115
timestamp 1667941163
transform 1 0 11684 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_157
timestamp 1667941163
transform 1 0 15548 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_178
timestamp 1667941163
transform 1 0 17480 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_186
timestamp 1667941163
transform 1 0 18216 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1667941163
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_205
timestamp 1667941163
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1667941163
transform 1 0 20424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1667941163
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1667941163
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1667941163
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_278
timestamp 1667941163
transform 1 0 26680 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_296
timestamp 1667941163
transform 1 0 28336 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_315
timestamp 1667941163
transform 1 0 30084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_323
timestamp 1667941163
transform 1 0 30820 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_328
timestamp 1667941163
transform 1 0 31280 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_335
timestamp 1667941163
transform 1 0 31924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_347
timestamp 1667941163
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1667941163
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_398
timestamp 1667941163
transform 1 0 37720 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_405
timestamp 1667941163
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_41
timestamp 1667941163
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_80
timestamp 1667941163
transform 1 0 8464 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_92
timestamp 1667941163
transform 1 0 9568 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1667941163
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_122
timestamp 1667941163
transform 1 0 12328 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_130
timestamp 1667941163
transform 1 0 13064 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_139
timestamp 1667941163
transform 1 0 13892 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_145
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1667941163
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1667941163
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_174
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_182
timestamp 1667941163
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_201
timestamp 1667941163
transform 1 0 19596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_213
timestamp 1667941163
transform 1 0 20700 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1667941163
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 1667941163
transform 1 0 23276 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_262
timestamp 1667941163
transform 1 0 25208 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_270
timestamp 1667941163
transform 1 0 25944 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1667941163
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_323
timestamp 1667941163
transform 1 0 30820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1667941163
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_400
timestamp 1667941163
transform 1 0 37904 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1667941163
transform 1 0 38456 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_38
timestamp 1667941163
transform 1 0 4600 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_48
timestamp 1667941163
transform 1 0 5520 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_60
timestamp 1667941163
transform 1 0 6624 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_72
timestamp 1667941163
transform 1 0 7728 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_91
timestamp 1667941163
transform 1 0 9476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_100
timestamp 1667941163
transform 1 0 10304 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_120
timestamp 1667941163
transform 1 0 12144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_127
timestamp 1667941163
transform 1 0 12788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_131
timestamp 1667941163
transform 1 0 13156 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_151
timestamp 1667941163
transform 1 0 14996 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_160
timestamp 1667941163
transform 1 0 15824 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_172
timestamp 1667941163
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_184
timestamp 1667941163
transform 1 0 18032 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_206
timestamp 1667941163
transform 1 0 20056 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_215
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_223
timestamp 1667941163
transform 1 0 21620 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_230
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_242
timestamp 1667941163
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1667941163
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_262
timestamp 1667941163
transform 1 0 25208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_274
timestamp 1667941163
transform 1 0 26312 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_279
timestamp 1667941163
transform 1 0 26772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_287
timestamp 1667941163
transform 1 0 27508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_295
timestamp 1667941163
transform 1 0 28244 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1667941163
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_314
timestamp 1667941163
transform 1 0 29992 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_328
timestamp 1667941163
transform 1 0 31280 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_336
timestamp 1667941163
transform 1 0 32016 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_342
timestamp 1667941163
transform 1 0 32568 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_354
timestamp 1667941163
transform 1 0 33672 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1667941163
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_383
timestamp 1667941163
transform 1 0 36340 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_14
timestamp 1667941163
transform 1 0 2392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_22
timestamp 1667941163
transform 1 0 3128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_30
timestamp 1667941163
transform 1 0 3864 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1667941163
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_77
timestamp 1667941163
transform 1 0 8188 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_88
timestamp 1667941163
transform 1 0 9200 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_96
timestamp 1667941163
transform 1 0 9936 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1667941163
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_121
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_129
timestamp 1667941163
transform 1 0 12972 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1667941163
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_179
timestamp 1667941163
transform 1 0 17572 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_188
timestamp 1667941163
transform 1 0 18400 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_196
timestamp 1667941163
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_204
timestamp 1667941163
transform 1 0 19872 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_218
timestamp 1667941163
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_234
timestamp 1667941163
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_241
timestamp 1667941163
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_252
timestamp 1667941163
transform 1 0 24288 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_264
timestamp 1667941163
transform 1 0 25392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1667941163
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_294
timestamp 1667941163
transform 1 0 28152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_314
timestamp 1667941163
transform 1 0 29992 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_326
timestamp 1667941163
transform 1 0 31096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_346
timestamp 1667941163
transform 1 0 32936 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_358
timestamp 1667941163
transform 1 0 34040 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_370
timestamp 1667941163
transform 1 0 35144 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_382
timestamp 1667941163
transform 1 0 36248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1667941163
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_399
timestamp 1667941163
transform 1 0 37812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1667941163
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_111
timestamp 1667941163
transform 1 0 11316 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_123
timestamp 1667941163
transform 1 0 12420 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_131
timestamp 1667941163
transform 1 0 13156 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_149
timestamp 1667941163
transform 1 0 14812 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_157
timestamp 1667941163
transform 1 0 15548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_178
timestamp 1667941163
transform 1 0 17480 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_186
timestamp 1667941163
transform 1 0 18216 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1667941163
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_203
timestamp 1667941163
transform 1 0 19780 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_215
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_227
timestamp 1667941163
transform 1 0 21988 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_232
timestamp 1667941163
transform 1 0 22448 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1667941163
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_285
timestamp 1667941163
transform 1 0 27324 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_291
timestamp 1667941163
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1667941163
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_317
timestamp 1667941163
transform 1 0 30268 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_329
timestamp 1667941163
transform 1 0 31372 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_341
timestamp 1667941163
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1667941163
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1667941163
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_383
timestamp 1667941163
transform 1 0 36340 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_14
timestamp 1667941163
transform 1 0 2392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_21
timestamp 1667941163
transform 1 0 3036 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_28
timestamp 1667941163
transform 1 0 3680 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_35
timestamp 1667941163
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_47
timestamp 1667941163
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_87
timestamp 1667941163
transform 1 0 9108 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_94
timestamp 1667941163
transform 1 0 9752 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_106
timestamp 1667941163
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_145
timestamp 1667941163
transform 1 0 14444 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1667941163
transform 1 0 15272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1667941163
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_189
timestamp 1667941163
transform 1 0 18492 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_201
timestamp 1667941163
transform 1 0 19596 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1667941163
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1667941163
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_263
timestamp 1667941163
transform 1 0 25300 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1667941163
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_291
timestamp 1667941163
transform 1 0 27876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_303
timestamp 1667941163
transform 1 0 28980 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_311
timestamp 1667941163
transform 1 0 29716 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_355
timestamp 1667941163
transform 1 0 33764 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_377
timestamp 1667941163
transform 1 0 35788 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1667941163
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_400
timestamp 1667941163
transform 1 0 37904 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1667941163
transform 1 0 38456 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_16
timestamp 1667941163
transform 1 0 2576 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_35
timestamp 1667941163
transform 1 0 4324 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_39
timestamp 1667941163
transform 1 0 4692 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_51
timestamp 1667941163
transform 1 0 5796 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_63
timestamp 1667941163
transform 1 0 6900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_75
timestamp 1667941163
transform 1 0 8004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_92
timestamp 1667941163
transform 1 0 9568 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_103
timestamp 1667941163
transform 1 0 10580 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_115
timestamp 1667941163
transform 1 0 11684 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_119
timestamp 1667941163
transform 1 0 12052 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1667941163
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_149
timestamp 1667941163
transform 1 0 14812 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_158
timestamp 1667941163
transform 1 0 15640 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_166
timestamp 1667941163
transform 1 0 16376 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_173
timestamp 1667941163
transform 1 0 17020 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_204
timestamp 1667941163
transform 1 0 19872 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_208
timestamp 1667941163
transform 1 0 20240 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_216
timestamp 1667941163
transform 1 0 20976 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_220
timestamp 1667941163
transform 1 0 21344 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_237
timestamp 1667941163
transform 1 0 22908 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1667941163
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_260
timestamp 1667941163
transform 1 0 25024 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_272
timestamp 1667941163
transform 1 0 26128 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_280
timestamp 1667941163
transform 1 0 26864 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_285
timestamp 1667941163
transform 1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1667941163
transform 1 0 28152 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_327
timestamp 1667941163
transform 1 0 31188 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_339
timestamp 1667941163
transform 1 0 32292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_351
timestamp 1667941163
transform 1 0 33396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_358
timestamp 1667941163
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1667941163
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_43
timestamp 1667941163
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_88
timestamp 1667941163
transform 1 0 9200 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1667941163
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_119
timestamp 1667941163
transform 1 0 12052 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_136
timestamp 1667941163
transform 1 0 13616 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_144
timestamp 1667941163
transform 1 0 14352 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_153
timestamp 1667941163
transform 1 0 15180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1667941163
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1667941163
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_190
timestamp 1667941163
transform 1 0 18584 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_196
timestamp 1667941163
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_211
timestamp 1667941163
transform 1 0 20516 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1667941163
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_255
timestamp 1667941163
transform 1 0 24564 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_264
timestamp 1667941163
transform 1 0 25392 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1667941163
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_289
timestamp 1667941163
transform 1 0 27692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_297
timestamp 1667941163
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_306
timestamp 1667941163
transform 1 0 29256 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_318
timestamp 1667941163
transform 1 0 30360 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_330
timestamp 1667941163
transform 1 0 31464 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_381
timestamp 1667941163
transform 1 0 36156 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1667941163
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_400
timestamp 1667941163
transform 1 0 37904 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1667941163
transform 1 0 38456 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_13
timestamp 1667941163
transform 1 0 2300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_25
timestamp 1667941163
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_104
timestamp 1667941163
transform 1 0 10672 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_116
timestamp 1667941163
transform 1 0 11776 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_124
timestamp 1667941163
transform 1 0 12512 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_129
timestamp 1667941163
transform 1 0 12972 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1667941163
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1667941163
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_164
timestamp 1667941163
transform 1 0 16192 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_181
timestamp 1667941163
transform 1 0 17756 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_212
timestamp 1667941163
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1667941163
transform 1 0 21620 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_227
timestamp 1667941163
transform 1 0 21988 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_232
timestamp 1667941163
transform 1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_240
timestamp 1667941163
transform 1 0 23184 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_262
timestamp 1667941163
transform 1 0 25208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_266
timestamp 1667941163
transform 1 0 25576 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_275
timestamp 1667941163
transform 1 0 26404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_287
timestamp 1667941163
transform 1 0 27508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_299
timestamp 1667941163
transform 1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_383
timestamp 1667941163
transform 1 0 36340 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_7
timestamp 1667941163
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_29
timestamp 1667941163
transform 1 0 3772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_41
timestamp 1667941163
transform 1 0 4876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1667941163
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_145
timestamp 1667941163
transform 1 0 14444 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_153
timestamp 1667941163
transform 1 0 15180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1667941163
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_177
timestamp 1667941163
transform 1 0 17388 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_189
timestamp 1667941163
transform 1 0 18492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_201
timestamp 1667941163
transform 1 0 19596 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_209
timestamp 1667941163
transform 1 0 20332 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1667941163
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_248
timestamp 1667941163
transform 1 0 23920 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_259
timestamp 1667941163
transform 1 0 24932 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_266
timestamp 1667941163
transform 1 0 25576 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1667941163
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_290
timestamp 1667941163
transform 1 0 27784 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_294
timestamp 1667941163
transform 1 0 28152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_306
timestamp 1667941163
transform 1 0 29256 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_318
timestamp 1667941163
transform 1 0 30360 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1667941163
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_342
timestamp 1667941163
transform 1 0 32568 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_350
timestamp 1667941163
transform 1 0 33304 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_374
timestamp 1667941163
transform 1 0 35512 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_383
timestamp 1667941163
transform 1 0 36340 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1667941163
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_398
timestamp 1667941163
transform 1 0 37720 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_12
timestamp 1667941163
transform 1 0 2208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1667941163
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_148
timestamp 1667941163
transform 1 0 14720 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_162
timestamp 1667941163
transform 1 0 16008 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_168
timestamp 1667941163
transform 1 0 16560 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1667941163
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_187
timestamp 1667941163
transform 1 0 18308 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1667941163
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_212
timestamp 1667941163
transform 1 0 20608 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_220
timestamp 1667941163
transform 1 0 21344 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_237
timestamp 1667941163
transform 1 0 22908 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_244
timestamp 1667941163
transform 1 0 23552 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_271
timestamp 1667941163
transform 1 0 26036 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_279
timestamp 1667941163
transform 1 0 26772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_286
timestamp 1667941163
transform 1 0 27416 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_293
timestamp 1667941163
transform 1 0 28060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1667941163
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_337
timestamp 1667941163
transform 1 0 32108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_359
timestamp 1667941163
transform 1 0 34132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_369
timestamp 1667941163
transform 1 0 35052 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_373
timestamp 1667941163
transform 1 0 35420 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_380
timestamp 1667941163
transform 1 0 36064 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_405
timestamp 1667941163
transform 1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_26
timestamp 1667941163
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_38
timestamp 1667941163
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1667941163
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_151
timestamp 1667941163
transform 1 0 14996 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_163
timestamp 1667941163
transform 1 0 16100 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_177
timestamp 1667941163
transform 1 0 17388 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_186
timestamp 1667941163
transform 1 0 18216 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_194
timestamp 1667941163
transform 1 0 18952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_208
timestamp 1667941163
transform 1 0 20240 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_240
timestamp 1667941163
transform 1 0 23184 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_265
timestamp 1667941163
transform 1 0 25484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1667941163
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_298
timestamp 1667941163
transform 1 0 28520 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_346
timestamp 1667941163
transform 1 0 32936 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_357
timestamp 1667941163
transform 1 0 33948 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1667941163
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_398
timestamp 1667941163
transform 1 0 37720 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_159
timestamp 1667941163
transform 1 0 15732 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_171
timestamp 1667941163
transform 1 0 16836 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_175
timestamp 1667941163
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_187
timestamp 1667941163
transform 1 0 18308 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1667941163
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_206
timestamp 1667941163
transform 1 0 20056 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1667941163
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_235
timestamp 1667941163
transform 1 0 22724 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_247
timestamp 1667941163
transform 1 0 23828 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_273
timestamp 1667941163
transform 1 0 26220 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_279
timestamp 1667941163
transform 1 0 26772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1667941163
transform 1 0 27416 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_290
timestamp 1667941163
transform 1 0 27784 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_294
timestamp 1667941163
transform 1 0 28152 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_313
timestamp 1667941163
transform 1 0 29900 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_317
timestamp 1667941163
transform 1 0 30268 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_324
timestamp 1667941163
transform 1 0 30912 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_335
timestamp 1667941163
transform 1 0 31924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_342
timestamp 1667941163
transform 1 0 32568 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_349
timestamp 1667941163
transform 1 0 33212 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1667941163
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_370
timestamp 1667941163
transform 1 0 35144 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_374
timestamp 1667941163
transform 1 0 35512 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_378
timestamp 1667941163
transform 1 0 35880 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_16
timestamp 1667941163
transform 1 0 2576 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_23
timestamp 1667941163
transform 1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_30
timestamp 1667941163
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_42
timestamp 1667941163
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1667941163
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_154
timestamp 1667941163
transform 1 0 15272 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_187
timestamp 1667941163
transform 1 0 18308 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_194
timestamp 1667941163
transform 1 0 18952 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_206
timestamp 1667941163
transform 1 0 20056 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_214
timestamp 1667941163
transform 1 0 20792 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1667941163
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1667941163
transform 1 0 23460 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_247
timestamp 1667941163
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_254
timestamp 1667941163
transform 1 0 24472 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_263
timestamp 1667941163
transform 1 0 25300 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_269
timestamp 1667941163
transform 1 0 25852 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_287
timestamp 1667941163
transform 1 0 27508 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_309
timestamp 1667941163
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_316
timestamp 1667941163
transform 1 0 30176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_323
timestamp 1667941163
transform 1 0 30820 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_330
timestamp 1667941163
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_343
timestamp 1667941163
transform 1 0 32660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_365
timestamp 1667941163
transform 1 0 34684 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_398
timestamp 1667941163
transform 1 0 37720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_52
timestamp 1667941163
transform 1 0 5888 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_56
timestamp 1667941163
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_60
timestamp 1667941163
transform 1 0 6624 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_72
timestamp 1667941163
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_92
timestamp 1667941163
transform 1 0 9568 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_104
timestamp 1667941163
transform 1 0 10672 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_116
timestamp 1667941163
transform 1 0 11776 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_128
timestamp 1667941163
transform 1 0 12880 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_147
timestamp 1667941163
transform 1 0 14628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_169
timestamp 1667941163
transform 1 0 16652 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1667941163
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_206
timestamp 1667941163
transform 1 0 20056 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_214
timestamp 1667941163
transform 1 0 20792 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1667941163
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_244
timestamp 1667941163
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_276
timestamp 1667941163
transform 1 0 26496 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_332
timestamp 1667941163
transform 1 0 31648 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_371
timestamp 1667941163
transform 1 0 35236 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_393
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_400
timestamp 1667941163
transform 1 0 37904 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1667941163
transform 1 0 38456 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_7
timestamp 1667941163
transform 1 0 1748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_29
timestamp 1667941163
transform 1 0 3772 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_80
timestamp 1667941163
transform 1 0 8464 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1667941163
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_175
timestamp 1667941163
transform 1 0 17204 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_197
timestamp 1667941163
transform 1 0 19228 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1667941163
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_304
timestamp 1667941163
transform 1 0 29072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_360
timestamp 1667941163
transform 1 0 34224 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1667941163
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_398
timestamp 1667941163
transform 1 0 37720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_16
timestamp 1667941163
transform 1 0 2576 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_22
timestamp 1667941163
transform 1 0 3128 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_74
timestamp 1667941163
transform 1 0 7912 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_91
timestamp 1667941163
transform 1 0 9476 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_103
timestamp 1667941163
transform 1 0 10580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1667941163
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_160
timestamp 1667941163
transform 1 0 15824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_180
timestamp 1667941163
transform 1 0 17664 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_187
timestamp 1667941163
transform 1 0 18308 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_214
timestamp 1667941163
transform 1 0 20792 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 1667941163
transform 1 0 21252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1667941163
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1667941163
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1667941163
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 3128 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4968 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0725_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 38088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 22080 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform -1 0 36984 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform -1 0 4876 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10304 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform -1 0 33212 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 37444 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 33672 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform -1 0 28428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 37444 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform -1 0 28152 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 26496 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0745_
timestamp 1667941163
transform 1 0 10028 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform -1 0 36984 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 37536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform -1 0 35144 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0752_
timestamp 1667941163
transform 1 0 4324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 2944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform -1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform -1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform -1 0 2300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform -1 0 3680 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0759_
timestamp 1667941163
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0760_
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform -1 0 17664 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform -1 0 2852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform -1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 23552 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform -1 0 15824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0767_
timestamp 1667941163
transform 1 0 2668 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 30544 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform -1 0 2576 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 38088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 37444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0774_
timestamp 1667941163
transform -1 0 4232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform -1 0 2576 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform -1 0 20056 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform -1 0 37720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform -1 0 2576 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 36432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform -1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 35880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0788_
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 23184 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform -1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0795_
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 35604 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 25944 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 37444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform -1 0 4600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 37444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform -1 0 36984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0802_
timestamp 1667941163
transform 1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0803_
timestamp 1667941163
transform -1 0 3496 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 23276 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 28520 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform -1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 25024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 9292 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform -1 0 15272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0810_
timestamp 1667941163
transform -1 0 4784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 20976 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 37444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform -1 0 2392 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0817_
timestamp 1667941163
transform 1 0 3772 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 6348 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 37444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform -1 0 2852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform -1 0 36340 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 37444 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0824_
timestamp 1667941163
transform 1 0 2852 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform -1 0 3128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform -1 0 30176 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 29992 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 33764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 33764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0831_
timestamp 1667941163
transform -1 0 4508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 32936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform -1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0838_
timestamp 1667941163
transform 1 0 5152 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 38088 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 31648 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform -1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 37444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform -1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0845_
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform -1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform -1 0 18952 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 32292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform -1 0 3220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform -1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform -1 0 2944 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20976 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform -1 0 20792 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22908 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 23276 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0858_
timestamp 1667941163
transform -1 0 21528 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0859_
timestamp 1667941163
transform 1 0 20240 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0860_
timestamp 1667941163
transform 1 0 22816 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19872 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0862_
timestamp 1667941163
transform 1 0 18584 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0864_
timestamp 1667941163
transform 1 0 18124 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19964 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 1667941163
transform 1 0 4416 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform -1 0 13064 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0869_
timestamp 1667941163
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0870_
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0871_
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0874_
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0875_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0876_
timestamp 1667941163
transform -1 0 13800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0877_
timestamp 1667941163
transform -1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0878_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18952 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0879_
timestamp 1667941163
transform -1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0880_
timestamp 1667941163
transform -1 0 13800 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18032 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0882_
timestamp 1667941163
transform -1 0 20976 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0883_
timestamp 1667941163
transform -1 0 14904 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0884_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11868 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0885_
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14168 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0887_
timestamp 1667941163
transform -1 0 20608 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0888_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0889_
timestamp 1667941163
transform 1 0 19044 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0890_
timestamp 1667941163
transform 1 0 20516 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1667941163
transform -1 0 35328 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0892_
timestamp 1667941163
transform -1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18032 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0894_
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12696 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18216 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0897_
timestamp 1667941163
transform -1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0898_
timestamp 1667941163
transform -1 0 9568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0899_
timestamp 1667941163
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0900_
timestamp 1667941163
transform 1 0 19228 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0901_
timestamp 1667941163
transform 1 0 16652 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20056 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0903_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19504 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0906_
timestamp 1667941163
transform 1 0 24840 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0907_
timestamp 1667941163
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26220 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1667941163
transform 1 0 25760 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0910_
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _0911_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0912_
timestamp 1667941163
transform 1 0 27140 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0913_
timestamp 1667941163
transform 1 0 26404 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1667941163
transform 1 0 29716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0915_
timestamp 1667941163
transform 1 0 29900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0916_
timestamp 1667941163
transform -1 0 28888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0917_
timestamp 1667941163
transform 1 0 27784 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0918_
timestamp 1667941163
transform 1 0 27140 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0919_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0920_
timestamp 1667941163
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1667941163
transform 1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14812 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0924_
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0925_
timestamp 1667941163
transform 1 0 15548 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0926_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0927_
timestamp 1667941163
transform 1 0 13340 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0928_
timestamp 1667941163
transform -1 0 15088 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0929_
timestamp 1667941163
transform 1 0 13156 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12788 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0932_
timestamp 1667941163
transform -1 0 13524 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0933_
timestamp 1667941163
transform 1 0 10580 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1667941163
transform 1 0 12512 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14996 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0936_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13432 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0937_
timestamp 1667941163
transform 1 0 8648 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0938_
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0939_
timestamp 1667941163
transform 1 0 9476 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0940_
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0941_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1667941163
transform -1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0945_
timestamp 1667941163
transform -1 0 8832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1667941163
transform -1 0 9476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0947_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0948_
timestamp 1667941163
transform 1 0 9292 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0949_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0950_
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0951_
timestamp 1667941163
transform 1 0 15088 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0953_
timestamp 1667941163
transform -1 0 15824 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0954_
timestamp 1667941163
transform -1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0955_
timestamp 1667941163
transform -1 0 9016 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0956_
timestamp 1667941163
transform -1 0 8188 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0957_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 8464 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0959_
timestamp 1667941163
transform 1 0 8004 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0960_
timestamp 1667941163
transform 1 0 8648 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0961_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14720 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0963_
timestamp 1667941163
transform -1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0964_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16008 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17296 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1667941163
transform 1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0967_
timestamp 1667941163
transform -1 0 17664 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0968_
timestamp 1667941163
transform 1 0 14996 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0969_
timestamp 1667941163
transform -1 0 17572 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0970_
timestamp 1667941163
transform 1 0 18584 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0971_
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0972_
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17296 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1667941163
transform 1 0 17940 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18216 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1667941163
transform -1 0 17296 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0977_
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0978_
timestamp 1667941163
transform 1 0 12696 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0979_
timestamp 1667941163
transform 1 0 13248 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0980_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 1667941163
transform 1 0 18032 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0982_
timestamp 1667941163
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0983_
timestamp 1667941163
transform 1 0 21160 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0984_
timestamp 1667941163
transform 1 0 18400 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0985_
timestamp 1667941163
transform -1 0 19964 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0986_
timestamp 1667941163
transform -1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0987_
timestamp 1667941163
transform -1 0 17664 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0988_
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17020 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform -1 0 18308 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0991_
timestamp 1667941163
transform 1 0 12420 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1667941163
transform 1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0993_
timestamp 1667941163
transform -1 0 13064 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 12696 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0995_
timestamp 1667941163
transform -1 0 12236 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0996_
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0997_
timestamp 1667941163
transform -1 0 12328 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform -1 0 10304 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0999_
timestamp 1667941163
transform 1 0 9936 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1000_
timestamp 1667941163
transform 1 0 10396 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1667941163
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1667941163
transform 1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1003_
timestamp 1667941163
transform -1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1004_
timestamp 1667941163
transform 1 0 16836 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1006_
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1667941163
transform -1 0 9660 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1008_
timestamp 1667941163
transform -1 0 20148 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1009_
timestamp 1667941163
transform -1 0 17848 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1010_
timestamp 1667941163
transform -1 0 10304 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1011_
timestamp 1667941163
transform 1 0 9384 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform -1 0 10488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1013_
timestamp 1667941163
transform -1 0 10304 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1667941163
transform -1 0 8648 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 9476 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1016_
timestamp 1667941163
transform -1 0 9568 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1018_
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1667941163
transform -1 0 9752 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1020_
timestamp 1667941163
transform 1 0 8740 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1021_
timestamp 1667941163
transform 1 0 8280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1022_
timestamp 1667941163
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1023_
timestamp 1667941163
transform 1 0 8740 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1024_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1025_
timestamp 1667941163
transform -1 0 10120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1026_
timestamp 1667941163
transform 1 0 9936 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1027_
timestamp 1667941163
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1028_
timestamp 1667941163
transform -1 0 10580 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1029_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1030_
timestamp 1667941163
transform 1 0 16008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1667941163
transform -1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1032_
timestamp 1667941163
transform 1 0 8740 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1667941163
transform -1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1034_
timestamp 1667941163
transform -1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1035_
timestamp 1667941163
transform 1 0 10212 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1036_
timestamp 1667941163
transform 1 0 12420 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1667941163
transform 1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1038_
timestamp 1667941163
transform -1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1039_
timestamp 1667941163
transform -1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1040_
timestamp 1667941163
transform 1 0 9384 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1041_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1042_
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1667941163
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1044_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1667941163
transform -1 0 17020 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1046_
timestamp 1667941163
transform 1 0 20976 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1047_
timestamp 1667941163
transform -1 0 18768 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1048_
timestamp 1667941163
transform -1 0 17572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1049_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1667941163
transform 1 0 17572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1667941163
transform -1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17020 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1667941163
transform -1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1667941163
transform 1 0 21160 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1057_
timestamp 1667941163
transform 1 0 14996 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1058_
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _1059_
timestamp 1667941163
transform -1 0 17848 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1061_
timestamp 1667941163
transform -1 0 12972 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1063_
timestamp 1667941163
transform 1 0 12788 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1064_
timestamp 1667941163
transform 1 0 10212 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1065_
timestamp 1667941163
transform 1 0 11224 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1066_
timestamp 1667941163
transform -1 0 14812 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1067_
timestamp 1667941163
transform -1 0 20240 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1068_
timestamp 1667941163
transform -1 0 14996 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1069_
timestamp 1667941163
transform -1 0 14720 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14628 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1071_
timestamp 1667941163
transform 1 0 14628 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1072_
timestamp 1667941163
transform -1 0 15640 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1073_
timestamp 1667941163
transform 1 0 15640 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1074_
timestamp 1667941163
transform -1 0 15272 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1667941163
transform 1 0 12696 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1076_
timestamp 1667941163
transform 1 0 20608 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1077_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1078_
timestamp 1667941163
transform -1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1079_
timestamp 1667941163
transform -1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1080_
timestamp 1667941163
transform -1 0 18492 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1081_
timestamp 1667941163
transform 1 0 18124 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1082_
timestamp 1667941163
transform -1 0 20332 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1083_
timestamp 1667941163
transform 1 0 20976 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1084_
timestamp 1667941163
transform 1 0 19964 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 1667941163
transform -1 0 21344 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1086_
timestamp 1667941163
transform 1 0 19412 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1087_
timestamp 1667941163
transform 1 0 20608 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1667941163
transform -1 0 20884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1089_
timestamp 1667941163
transform -1 0 18952 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1090_
timestamp 1667941163
transform 1 0 18400 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1091_
timestamp 1667941163
transform -1 0 18216 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1667941163
transform 1 0 16928 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1093_
timestamp 1667941163
transform 1 0 16836 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1094_
timestamp 1667941163
transform 1 0 16652 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1095_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1096_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1097_
timestamp 1667941163
transform 1 0 22080 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1098_
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1099_
timestamp 1667941163
transform -1 0 25208 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1100_
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1101_
timestamp 1667941163
transform -1 0 19872 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1102_
timestamp 1667941163
transform -1 0 19044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1103_
timestamp 1667941163
transform 1 0 26404 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1667941163
transform -1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1106_
timestamp 1667941163
transform 1 0 18952 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1107_
timestamp 1667941163
transform 1 0 22448 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1108_
timestamp 1667941163
transform 1 0 19228 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1109_
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1110_
timestamp 1667941163
transform 1 0 20516 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1111_
timestamp 1667941163
transform -1 0 26220 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1112_
timestamp 1667941163
transform -1 0 25392 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1113_
timestamp 1667941163
transform -1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1114_
timestamp 1667941163
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1115_
timestamp 1667941163
transform -1 0 24104 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1116_
timestamp 1667941163
transform -1 0 22540 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1117_
timestamp 1667941163
transform 1 0 23920 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1119_
timestamp 1667941163
transform -1 0 24564 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23736 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1121_
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1122_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20148 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1123_
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1667941163
transform 1 0 21252 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1125_
timestamp 1667941163
transform -1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1667941163
transform 1 0 20976 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1127_
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1128_
timestamp 1667941163
transform -1 0 21436 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1129_
timestamp 1667941163
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1130_
timestamp 1667941163
transform 1 0 30544 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1131_
timestamp 1667941163
transform -1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1667941163
transform -1 0 21436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1133_
timestamp 1667941163
transform -1 0 20976 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1134_
timestamp 1667941163
transform -1 0 24104 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1135_
timestamp 1667941163
transform -1 0 23276 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1136_
timestamp 1667941163
transform -1 0 22264 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1137_
timestamp 1667941163
transform -1 0 22632 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1138_
timestamp 1667941163
transform -1 0 22448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 1667941163
transform -1 0 27416 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1140_
timestamp 1667941163
transform 1 0 26956 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1141_
timestamp 1667941163
transform -1 0 28060 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1142_
timestamp 1667941163
transform 1 0 27232 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1143_
timestamp 1667941163
transform -1 0 29256 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1144_
timestamp 1667941163
transform 1 0 25760 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1145_
timestamp 1667941163
transform -1 0 28152 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1146_
timestamp 1667941163
transform 1 0 23276 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1147_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1148_
timestamp 1667941163
transform 1 0 23644 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1149_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1151_
timestamp 1667941163
transform 1 0 27232 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1152_
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1153_
timestamp 1667941163
transform -1 0 28888 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1154_
timestamp 1667941163
transform 1 0 25668 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1155_
timestamp 1667941163
transform 1 0 26772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1156_
timestamp 1667941163
transform -1 0 27876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1157_
timestamp 1667941163
transform -1 0 28152 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1158_
timestamp 1667941163
transform -1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1159_
timestamp 1667941163
transform 1 0 27876 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27140 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1162_
timestamp 1667941163
transform 1 0 28520 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1667941163
transform 1 0 24380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1164_
timestamp 1667941163
transform 1 0 25576 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1667941163
transform -1 0 25300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1166_
timestamp 1667941163
transform -1 0 25208 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1167_
timestamp 1667941163
transform 1 0 25668 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 1667941163
transform 1 0 24472 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1667941163
transform -1 0 25576 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1170_
timestamp 1667941163
transform -1 0 24012 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1171_
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1172_
timestamp 1667941163
transform 1 0 20608 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1667941163
transform -1 0 21528 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1174_
timestamp 1667941163
transform 1 0 14536 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1175_
timestamp 1667941163
transform 1 0 15548 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _1176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17940 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1177_
timestamp 1667941163
transform 1 0 23460 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1178_
timestamp 1667941163
transform -1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1179_
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1667941163
transform 1 0 28980 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1181_
timestamp 1667941163
transform 1 0 29808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1182_
timestamp 1667941163
transform -1 0 24564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1667941163
transform 1 0 17756 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1184_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1667941163
transform 1 0 22724 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1667941163
transform -1 0 24656 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 1667941163
transform 1 0 22816 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1188_
timestamp 1667941163
transform -1 0 23828 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1189_
timestamp 1667941163
transform 1 0 23460 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1190_
timestamp 1667941163
transform 1 0 23460 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1191_
timestamp 1667941163
transform -1 0 24932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1192_
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1193_
timestamp 1667941163
transform 1 0 31188 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1667941163
transform -1 0 32752 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1195_
timestamp 1667941163
transform 1 0 32200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1667941163
transform -1 0 32568 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1197_
timestamp 1667941163
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1198_
timestamp 1667941163
transform 1 0 30544 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1199_
timestamp 1667941163
transform -1 0 30268 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1667941163
transform 1 0 31648 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1201_
timestamp 1667941163
transform 1 0 30912 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1202_
timestamp 1667941163
transform 1 0 30360 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1203_
timestamp 1667941163
transform 1 0 30544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1204_
timestamp 1667941163
transform 1 0 31188 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1205_
timestamp 1667941163
transform -1 0 31832 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1206_
timestamp 1667941163
transform -1 0 32936 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1207_
timestamp 1667941163
transform 1 0 30360 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1208_
timestamp 1667941163
transform -1 0 29992 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1209_
timestamp 1667941163
transform 1 0 29808 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1210_
timestamp 1667941163
transform 1 0 30084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1211_
timestamp 1667941163
transform -1 0 31464 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1212_
timestamp 1667941163
transform 1 0 30544 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1213_
timestamp 1667941163
transform 1 0 31280 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1214_
timestamp 1667941163
transform 1 0 30912 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1215_
timestamp 1667941163
transform 1 0 29808 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1216_
timestamp 1667941163
transform 1 0 28980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp 1667941163
transform 1 0 28152 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1218_
timestamp 1667941163
transform 1 0 29716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1219_
timestamp 1667941163
transform -1 0 29348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1667941163
transform -1 0 29624 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1222_
timestamp 1667941163
transform -1 0 28980 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1223_
timestamp 1667941163
transform -1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1224_
timestamp 1667941163
transform 1 0 24656 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1225_
timestamp 1667941163
transform 1 0 30544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1227_
timestamp 1667941163
transform 1 0 26220 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1228_
timestamp 1667941163
transform -1 0 26680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1229_
timestamp 1667941163
transform -1 0 26956 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1230_
timestamp 1667941163
transform -1 0 25944 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1231_
timestamp 1667941163
transform 1 0 24656 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1232_
timestamp 1667941163
transform 1 0 25116 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1234_
timestamp 1667941163
transform -1 0 26404 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1235_
timestamp 1667941163
transform -1 0 27048 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1236_
timestamp 1667941163
transform -1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1237_
timestamp 1667941163
transform -1 0 26220 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1238_
timestamp 1667941163
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1239_
timestamp 1667941163
transform -1 0 21528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1240_
timestamp 1667941163
transform 1 0 26404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27416 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1242_
timestamp 1667941163
transform -1 0 27600 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1243_
timestamp 1667941163
transform 1 0 30452 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1244_
timestamp 1667941163
transform -1 0 32108 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1245_
timestamp 1667941163
transform 1 0 30360 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1246_
timestamp 1667941163
transform -1 0 29808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1247_
timestamp 1667941163
transform -1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1248_
timestamp 1667941163
transform -1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1249_
timestamp 1667941163
transform -1 0 15088 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1250_
timestamp 1667941163
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _1251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17756 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1252_
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17572 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1667941163
transform -1 0 22356 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1255_
timestamp 1667941163
transform -1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1256_
timestamp 1667941163
transform -1 0 18032 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1257_
timestamp 1667941163
transform -1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1258_
timestamp 1667941163
transform 1 0 17848 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1259_
timestamp 1667941163
transform 1 0 13800 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1260_
timestamp 1667941163
transform -1 0 14628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1261_
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1262_
timestamp 1667941163
transform -1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1263_
timestamp 1667941163
transform 1 0 17940 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1264_
timestamp 1667941163
transform -1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1265_
timestamp 1667941163
transform -1 0 16376 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1266_
timestamp 1667941163
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1267_
timestamp 1667941163
transform -1 0 19136 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1268_
timestamp 1667941163
transform -1 0 20424 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1269_
timestamp 1667941163
transform -1 0 20332 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1270_
timestamp 1667941163
transform -1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1271_
timestamp 1667941163
transform -1 0 20516 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1272_
timestamp 1667941163
transform 1 0 19872 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 1667941163
transform -1 0 19504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1667941163
transform -1 0 23000 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1275_
timestamp 1667941163
transform 1 0 20240 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1276_
timestamp 1667941163
transform -1 0 22448 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1277_
timestamp 1667941163
transform -1 0 21528 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1278_
timestamp 1667941163
transform 1 0 21712 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1279_
timestamp 1667941163
transform -1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1280_
timestamp 1667941163
transform 1 0 19504 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1281_
timestamp 1667941163
transform -1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1282_
timestamp 1667941163
transform -1 0 17480 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1283_
timestamp 1667941163
transform -1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1284_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1285_
timestamp 1667941163
transform -1 0 16376 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1286_
timestamp 1667941163
transform -1 0 16652 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1287_
timestamp 1667941163
transform -1 0 17480 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1288_
timestamp 1667941163
transform -1 0 16100 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1289_
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1290_
timestamp 1667941163
transform -1 0 15180 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1292_
timestamp 1667941163
transform -1 0 12788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1293_
timestamp 1667941163
transform 1 0 8924 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1667941163
transform 1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1667941163
transform -1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1296_
timestamp 1667941163
transform 1 0 11776 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1297_
timestamp 1667941163
transform -1 0 12144 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1667941163
transform -1 0 10672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1299_
timestamp 1667941163
transform 1 0 10212 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1300_
timestamp 1667941163
transform -1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1301_
timestamp 1667941163
transform -1 0 13340 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1302_
timestamp 1667941163
transform -1 0 13064 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1667941163
transform -1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14168 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 1667941163
transform 1 0 14076 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1306_
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1307_
timestamp 1667941163
transform -1 0 24472 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1308_
timestamp 1667941163
transform -1 0 28704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1667941163
transform -1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1667941163
transform 1 0 26036 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1311_
timestamp 1667941163
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 1667941163
transform -1 0 27600 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1313_
timestamp 1667941163
transform 1 0 26956 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1314_
timestamp 1667941163
transform -1 0 28060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1315_
timestamp 1667941163
transform -1 0 27692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1316_
timestamp 1667941163
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1317_
timestamp 1667941163
transform 1 0 30728 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1318_
timestamp 1667941163
transform 1 0 31556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1319_
timestamp 1667941163
transform 1 0 32292 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1320_
timestamp 1667941163
transform -1 0 28612 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1321_
timestamp 1667941163
transform 1 0 28060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1322_
timestamp 1667941163
transform 1 0 27232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1323_
timestamp 1667941163
transform 1 0 30544 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1324_
timestamp 1667941163
transform 1 0 31464 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1325_
timestamp 1667941163
transform -1 0 31832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1326_
timestamp 1667941163
transform 1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1327_
timestamp 1667941163
transform -1 0 32200 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1328_
timestamp 1667941163
transform 1 0 30360 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1667941163
transform -1 0 29992 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1330_
timestamp 1667941163
transform -1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1331_
timestamp 1667941163
transform 1 0 30544 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1332_
timestamp 1667941163
transform 1 0 30176 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1333_
timestamp 1667941163
transform -1 0 30728 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 1667941163
transform 1 0 31096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1335_
timestamp 1667941163
transform 1 0 30084 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1336_
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1337_
timestamp 1667941163
transform -1 0 29256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1338_
timestamp 1667941163
transform 1 0 27140 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1667941163
transform -1 0 31372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1340_
timestamp 1667941163
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1341_
timestamp 1667941163
transform -1 0 28520 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1342_
timestamp 1667941163
transform 1 0 26864 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1667941163
transform -1 0 22356 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1344_
timestamp 1667941163
transform 1 0 22724 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1345_
timestamp 1667941163
transform 1 0 27324 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1346_
timestamp 1667941163
transform -1 0 28796 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1667941163
transform -1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1348_
timestamp 1667941163
transform -1 0 28336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1349_
timestamp 1667941163
transform 1 0 28704 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1350_
timestamp 1667941163
transform -1 0 28520 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1351_
timestamp 1667941163
transform 1 0 27232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1352_
timestamp 1667941163
transform -1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1667941163
transform 1 0 27600 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1354_
timestamp 1667941163
transform 1 0 24932 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1355_
timestamp 1667941163
transform 1 0 25944 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1356_
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1357_
timestamp 1667941163
transform -1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20976 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1667941163
transform -1 0 18492 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1667941163
transform 1 0 12420 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1667941163
transform 1 0 10672 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1667941163
transform -1 0 11224 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1667941163
transform -1 0 19780 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1667941163
transform 1 0 14720 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1667941163
transform 1 0 10304 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1366_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10764 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1369_
timestamp 1667941163
transform 1 0 11684 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1667941163
transform 1 0 12144 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1667941163
transform 1 0 10764 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1667941163
transform 1 0 10672 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1667941163
transform 1 0 13800 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1667941163
transform 1 0 14352 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1667941163
transform 1 0 12144 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1667941163
transform -1 0 13616 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1378_
timestamp 1667941163
transform 1 0 18032 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1667941163
transform 1 0 21252 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1667941163
transform -1 0 21528 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1667941163
transform -1 0 26036 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1667941163
transform 1 0 22356 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1667941163
transform 1 0 21160 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1667941163
transform 1 0 29716 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1667941163
transform -1 0 29992 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1667941163
transform 1 0 28704 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1667941163
transform 1 0 27876 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1667941163
transform 1 0 24472 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1667941163
transform 1 0 25208 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1397_
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1667941163
transform 1 0 17848 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1667941163
transform -1 0 21160 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1667941163
transform -1 0 23552 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1667941163
transform 1 0 14904 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1667941163
transform 1 0 10304 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1667941163
transform 1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1667941163
transform -1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1667941163
transform 1 0 27692 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1667941163
transform 1 0 28704 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1667941163
transform -1 0 26772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1667941163
transform 1 0 22172 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1667941163
transform -1 0 25024 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1414_
timestamp 1667941163
transform 1 0 24380 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _1510__11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 2392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2116 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1511_
timestamp 1667941163
transform 1 0 1840 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1511__12
timestamp 1667941163
transform -1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1512__13
timestamp 1667941163
transform -1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1512_
timestamp 1667941163
transform 1 0 27876 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1513__14
timestamp 1667941163
transform 1 0 37628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1513_
timestamp 1667941163
transform -1 0 38364 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1514__15
timestamp 1667941163
transform -1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1514_
timestamp 1667941163
transform 1 0 8188 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1515__16
timestamp 1667941163
transform -1 0 13248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1515_
timestamp 1667941163
transform 1 0 12880 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1516__17
timestamp 1667941163
transform -1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1516_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1517__18
timestamp 1667941163
transform -1 0 37812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1517_
timestamp 1667941163
transform 1 0 36432 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1518__19
timestamp 1667941163
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1518_
timestamp 1667941163
transform 1 0 24288 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1519__20
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1519_
timestamp 1667941163
transform -1 0 29532 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1520_
timestamp 1667941163
transform 1 0 26864 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1520__21
timestamp 1667941163
transform -1 0 27416 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1521__22
timestamp 1667941163
transform -1 0 37904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1521_
timestamp 1667941163
transform 1 0 36432 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1522__23
timestamp 1667941163
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1522_
timestamp 1667941163
transform 1 0 8832 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1523__24
timestamp 1667941163
transform 1 0 37628 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1523_
timestamp 1667941163
transform -1 0 38364 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1524__25
timestamp 1667941163
transform -1 0 37720 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1524_
timestamp 1667941163
transform -1 0 37260 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1525__26
timestamp 1667941163
transform 1 0 36708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1525_
timestamp 1667941163
transform -1 0 36984 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1526_
timestamp 1667941163
transform 1 0 34592 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1526__27
timestamp 1667941163
transform 1 0 34132 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1527_
timestamp 1667941163
transform -1 0 3496 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1527__28
timestamp 1667941163
transform 1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1528__29
timestamp 1667941163
transform 1 0 2760 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1667941163
transform -1 0 3772 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1529__30
timestamp 1667941163
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1667941163
transform 1 0 5520 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1530__31
timestamp 1667941163
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1667941163
transform 1 0 1840 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1531__32
timestamp 1667941163
transform -1 0 2208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1532__33
timestamp 1667941163
transform 1 0 2024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1667941163
transform -1 0 3956 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1533__34
timestamp 1667941163
transform 1 0 18676 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1667941163
transform -1 0 18952 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1667941163
transform -1 0 3864 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1534__35
timestamp 1667941163
transform 1 0 3220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1535__36
timestamp 1667941163
transform -1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1536__37
timestamp 1667941163
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1667941163
transform 1 0 24564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1537__38
timestamp 1667941163
transform 1 0 24196 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1538__39
timestamp 1667941163
transform -1 0 15180 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1667941163
transform 1 0 14444 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1539__40
timestamp 1667941163
transform -1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1667941163
transform 1 0 19504 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1667941163
transform 1 0 32016 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1540__41
timestamp 1667941163
transform 1 0 31188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1541__42
timestamp 1667941163
transform -1 0 1932 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1667941163
transform -1 0 38364 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1542__43
timestamp 1667941163
transform 1 0 37628 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1543__44
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1667941163
transform -1 0 3772 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1544__45
timestamp 1667941163
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1667941163
transform -1 0 4048 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1545__46
timestamp 1667941163
transform 1 0 37628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1667941163
transform -1 0 38364 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1546__47
timestamp 1667941163
transform -1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1667941163
transform 1 0 5336 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1547__48
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1548__49
timestamp 1667941163
transform -1 0 20056 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1667941163
transform 1 0 19596 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1549__50
timestamp 1667941163
transform -1 0 37720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1667941163
transform 1 0 36432 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1550__51
timestamp 1667941163
transform 1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1667941163
transform -1 0 38364 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1551__52
timestamp 1667941163
transform -1 0 1932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1552__53
timestamp 1667941163
transform -1 0 37720 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1667941163
transform 1 0 36432 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1553__54
timestamp 1667941163
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1667941163
transform -1 0 3772 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1554__55
timestamp 1667941163
transform -1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1667941163
transform 1 0 20700 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1555_
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1555__56
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1556_
timestamp 1667941163
transform 1 0 23552 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1557_
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1558_
timestamp 1667941163
transform 1 0 3956 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1559_
timestamp 1667941163
transform 1 0 3864 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1560_
timestamp 1667941163
transform 1 0 14168 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1561_
timestamp 1667941163
transform 1 0 23828 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1562_
timestamp 1667941163
transform 1 0 33580 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1563_
timestamp 1667941163
transform -1 0 3496 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1564__57
timestamp 1667941163
transform -1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1564_
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1565__58
timestamp 1667941163
transform -1 0 37720 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1565_
timestamp 1667941163
transform -1 0 36984 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1566__59
timestamp 1667941163
transform -1 0 28060 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1566_
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1567__60
timestamp 1667941163
transform 1 0 38088 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1567_
timestamp 1667941163
transform -1 0 38364 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1568__61
timestamp 1667941163
transform -1 0 4324 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1568_
timestamp 1667941163
transform 1 0 4048 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1667941163
transform -1 0 38364 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1569__62
timestamp 1667941163
transform 1 0 37628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1570__63
timestamp 1667941163
transform -1 0 38364 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1667941163
transform 1 0 36432 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1571__64
timestamp 1667941163
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1667941163
transform 1 0 24380 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1572_
timestamp 1667941163
transform 1 0 29440 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1572__65
timestamp 1667941163
transform 1 0 28244 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1573_
timestamp 1667941163
transform -1 0 3496 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1573__66
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1574__67
timestamp 1667941163
transform -1 0 27416 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1574_
timestamp 1667941163
transform -1 0 26680 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1575__68
timestamp 1667941163
transform -1 0 9476 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1575_
timestamp 1667941163
transform 1 0 9200 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1576__69
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1576_
timestamp 1667941163
transform 1 0 14720 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1577__70
timestamp 1667941163
transform -1 0 21252 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1577_
timestamp 1667941163
transform 1 0 20976 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1578_
timestamp 1667941163
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1578__71
timestamp 1667941163
transform -1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1579__72
timestamp 1667941163
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1667941163
transform -1 0 3496 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1580__73
timestamp 1667941163
transform -1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1580_
timestamp 1667941163
transform -1 0 36984 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1581__74
timestamp 1667941163
transform -1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1581_
timestamp 1667941163
transform 1 0 25852 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1582_
timestamp 1667941163
transform -1 0 38272 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1582__75
timestamp 1667941163
transform -1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1583__76
timestamp 1667941163
transform 1 0 2760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1583_
timestamp 1667941163
transform -1 0 3496 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1584__77
timestamp 1667941163
transform -1 0 6808 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1584_
timestamp 1667941163
transform 1 0 6532 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1585__78
timestamp 1667941163
transform 1 0 38088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1585_
timestamp 1667941163
transform -1 0 38364 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1586__79
timestamp 1667941163
transform -1 0 2208 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1586_
timestamp 1667941163
transform 1 0 1840 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1587__80
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1587_
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1588_
timestamp 1667941163
transform -1 0 34684 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1588__81
timestamp 1667941163
transform -1 0 35420 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1589__82
timestamp 1667941163
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1589_
timestamp 1667941163
transform -1 0 38364 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1590__83
timestamp 1667941163
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1590_
timestamp 1667941163
transform -1 0 3772 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1591_
timestamp 1667941163
transform 1 0 29716 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1591__84
timestamp 1667941163
transform 1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1592__85
timestamp 1667941163
transform -1 0 34224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1592_
timestamp 1667941163
transform 1 0 33948 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1593_
timestamp 1667941163
transform 1 0 29900 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1593__86
timestamp 1667941163
transform -1 0 30912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1594_
timestamp 1667941163
transform 1 0 33856 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1595_
timestamp 1667941163
transform 1 0 33856 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1596_
timestamp 1667941163
transform 1 0 33580 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1597_
timestamp 1667941163
transform -1 0 11868 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1598_
timestamp 1667941163
transform 1 0 18400 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1599_
timestamp 1667941163
transform 1 0 32200 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1600__87
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1600_
timestamp 1667941163
transform -1 0 3496 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1601__88
timestamp 1667941163
transform -1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1601_
timestamp 1667941163
transform -1 0 3496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1602__89
timestamp 1667941163
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1602_
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1603_
timestamp 1667941163
transform -1 0 36984 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1603__90
timestamp 1667941163
transform -1 0 37904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1604_
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1604__91
timestamp 1667941163
transform -1 0 32568 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1605__92
timestamp 1667941163
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1605_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1606__93
timestamp 1667941163
transform -1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1606_
timestamp 1667941163
transform 1 0 11776 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1607__94
timestamp 1667941163
transform 1 0 37628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1607_
timestamp 1667941163
transform -1 0 38364 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1608__95
timestamp 1667941163
transform -1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1608_
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1609_
timestamp 1667941163
transform 1 0 1564 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1609__96
timestamp 1667941163
transform -1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1610__97
timestamp 1667941163
transform 1 0 18032 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1610_
timestamp 1667941163
transform -1 0 19228 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1611__98
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1611_
timestamp 1667941163
transform 1 0 4140 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1612_
timestamp 1667941163
transform -1 0 36984 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1612__99
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1613__100
timestamp 1667941163
transform -1 0 23000 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1613_
timestamp 1667941163
transform 1 0 22080 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1614_
timestamp 1667941163
transform 1 0 36432 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1614__101
timestamp 1667941163
transform -1 0 38364 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1615__102
timestamp 1667941163
transform 1 0 38088 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1615_
timestamp 1667941163
transform -1 0 38364 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1616_
timestamp 1667941163
transform 1 0 4232 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1616__103
timestamp 1667941163
transform -1 0 4600 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1617_
timestamp 1667941163
transform 1 0 32476 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1617__104
timestamp 1667941163
transform -1 0 32936 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1618__105
timestamp 1667941163
transform 1 0 38088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1618_
timestamp 1667941163
transform -1 0 38364 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1667941163
transform -1 0 17480 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1667941163
transform -1 0 14812 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1667941163
transform -1 0 22632 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1667941163
transform 1 0 15640 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1667941163
transform -1 0 17480 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1667941163
transform 1 0 23368 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp 1667941163
transform -1 0 30084 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout9
timestamp 1667941163
transform 1 0 29532 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout10
timestamp 1667941163
transform -1 0 21252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform -1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform -1 0 38364 0 1 36992
box -38 -48 958 592
<< labels >>
flabel metal2 s -10 39200 102 39800 0 FreeSans 448 90 0 0 active
port 0 nsew signal input
flabel metal3 s 39200 11508 39800 11748 0 FreeSans 960 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 30902 200 31014 800 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal3 s 39200 6068 39800 6308 0 FreeSans 960 0 0 0 io_in[13]
port 5 nsew signal input
flabel metal3 s 39200 4028 39800 4268 0 FreeSans 960 0 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 200 5388 800 5628 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal3 s 39200 19668 39800 19908 0 FreeSans 960 0 0 0 io_in[17]
port 9 nsew signal input
flabel metal3 s 39200 14908 39800 15148 0 FreeSans 960 0 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 32190 200 32302 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 12226 39200 12338 39800 0 FreeSans 448 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 39200 628 39800 868 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 39200 29188 39800 29428 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 5142 39200 5254 39800 0 FreeSans 448 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 33478 39200 33590 39800 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal3 s 200 27148 800 27388 0 FreeSans 960 0 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 36698 39200 36810 39800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 18666 39200 18778 39800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 30258 200 30370 800 0 FreeSans 448 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 25750 200 25862 800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 7718 39200 7830 39800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 1278 39200 1390 39800 0 FreeSans 448 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 10294 39200 10406 39800 0 FreeSans 448 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal3 s 200 16268 800 16508 0 FreeSans 960 0 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 39200 1308 39800 1548 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 20598 200 20710 800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal3 s 39200 13548 39800 13788 0 FreeSans 960 0 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal3 s 39200 26468 39800 26708 0 FreeSans 960 0 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 33478 200 33590 800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 200 32588 800 32828 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 32834 200 32946 800 0 FreeSans 448 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal bidirectional
flabel metal2 s 28970 39200 29082 39800 0 FreeSans 448 90 0 0 io_oeb[10]
port 40 nsew signal bidirectional
flabel metal2 s 34766 200 34878 800 0 FreeSans 448 90 0 0 io_oeb[11]
port 41 nsew signal bidirectional
flabel metal2 s 30258 39200 30370 39800 0 FreeSans 448 90 0 0 io_oeb[12]
port 42 nsew signal bidirectional
flabel metal3 s 39200 23748 39800 23988 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal bidirectional
flabel metal3 s 39200 31908 39800 32148 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal bidirectional
flabel metal3 s 39200 23068 39800 23308 0 FreeSans 960 0 0 0 io_oeb[15]
port 45 nsew signal bidirectional
flabel metal3 s 200 12868 800 13108 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal bidirectional
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal bidirectional
flabel metal2 s 35410 39200 35522 39800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal bidirectional
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 io_oeb[19]
port 49 nsew signal bidirectional
flabel metal3 s 39200 1988 39800 2228 0 FreeSans 960 0 0 0 io_oeb[1]
port 50 nsew signal bidirectional
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal bidirectional
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal bidirectional
flabel metal3 s 39200 36668 39800 36908 0 FreeSans 960 0 0 0 io_oeb[22]
port 53 nsew signal bidirectional
flabel metal2 s 32190 39200 32302 39800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal bidirectional
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal bidirectional
flabel metal2 s 12226 200 12338 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal bidirectional
flabel metal3 s 39200 22388 39800 22628 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal bidirectional
flabel metal2 s 25106 200 25218 800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal bidirectional
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 io_oeb[28]
port 59 nsew signal bidirectional
flabel metal2 s 18022 39200 18134 39800 0 FreeSans 448 90 0 0 io_oeb[29]
port 60 nsew signal bidirectional
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 io_oeb[2]
port 61 nsew signal bidirectional
flabel metal2 s 3210 39200 3322 39800 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal bidirectional
flabel metal2 s 38630 39200 38742 39800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal bidirectional
flabel metal2 s 22530 39200 22642 39800 0 FreeSans 448 90 0 0 io_oeb[32]
port 64 nsew signal bidirectional
flabel metal3 s 39200 33948 39800 34188 0 FreeSans 960 0 0 0 io_oeb[33]
port 65 nsew signal bidirectional
flabel metal3 s 39200 34628 39800 34868 0 FreeSans 960 0 0 0 io_oeb[34]
port 66 nsew signal bidirectional
flabel metal3 s 200 19668 800 19908 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal bidirectional
flabel metal2 s 32834 39200 32946 39800 0 FreeSans 448 90 0 0 io_oeb[36]
port 68 nsew signal bidirectional
flabel metal3 s 39200 25108 39800 25348 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal bidirectional
flabel metal2 s 7074 39200 7186 39800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal bidirectional
flabel metal3 s 39200 10828 39800 11068 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal bidirectional
flabel metal3 s 200 33268 800 33508 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal bidirectional
flabel metal2 s 3854 39200 3966 39800 0 FreeSans 448 90 0 0 io_oeb[6]
port 73 nsew signal bidirectional
flabel metal3 s 39200 37348 39800 37588 0 FreeSans 960 0 0 0 io_oeb[7]
port 74 nsew signal bidirectional
flabel metal3 s 39200 18988 39800 19228 0 FreeSans 960 0 0 0 io_oeb[8]
port 75 nsew signal bidirectional
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[9]
port 76 nsew signal bidirectional
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal bidirectional
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal bidirectional
flabel metal2 s 21242 200 21354 800 0 FreeSans 448 90 0 0 io_out[11]
port 79 nsew signal bidirectional
flabel metal3 s 200 17628 800 17868 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal bidirectional
flabel metal2 s 24462 39200 24574 39800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal bidirectional
flabel metal2 s 39274 39200 39386 39800 0 FreeSans 448 90 0 0 io_out[14]
port 82 nsew signal bidirectional
flabel metal3 s 200 26468 800 26708 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal bidirectional
flabel metal2 s 3854 200 3966 800 0 FreeSans 448 90 0 0 io_out[16]
port 84 nsew signal bidirectional
flabel metal2 s 14802 39200 14914 39800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal bidirectional
flabel metal3 s 39200 8788 39800 9028 0 FreeSans 960 0 0 0 io_out[18]
port 86 nsew signal bidirectional
flabel metal2 s 34122 39200 34234 39800 0 FreeSans 448 90 0 0 io_out[19]
port 87 nsew signal bidirectional
flabel metal3 s 200 1988 800 2228 0 FreeSans 960 0 0 0 io_out[1]
port 88 nsew signal bidirectional
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_out[20]
port 89 nsew signal bidirectional
flabel metal2 s 34122 200 34234 800 0 FreeSans 448 90 0 0 io_out[21]
port 90 nsew signal bidirectional
flabel metal2 s 37986 39200 38098 39800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal bidirectional
flabel metal2 s 26394 39200 26506 39800 0 FreeSans 448 90 0 0 io_out[23]
port 92 nsew signal bidirectional
flabel metal3 s 39200 24428 39800 24668 0 FreeSans 960 0 0 0 io_out[24]
port 93 nsew signal bidirectional
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 io_out[25]
port 94 nsew signal bidirectional
flabel metal2 s 39274 200 39386 800 0 FreeSans 448 90 0 0 io_out[26]
port 95 nsew signal bidirectional
flabel metal3 s 39200 16948 39800 17188 0 FreeSans 960 0 0 0 io_out[27]
port 96 nsew signal bidirectional
flabel metal2 s 23818 39200 23930 39800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal bidirectional
flabel metal2 s 29614 39200 29726 39800 0 FreeSans 448 90 0 0 io_out[29]
port 98 nsew signal bidirectional
flabel metal3 s 39200 12868 39800 13108 0 FreeSans 960 0 0 0 io_out[2]
port 99 nsew signal bidirectional
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal bidirectional
flabel metal2 s 25750 39200 25862 39800 0 FreeSans 448 90 0 0 io_out[31]
port 101 nsew signal bidirectional
flabel metal2 s 9650 39200 9762 39800 0 FreeSans 448 90 0 0 io_out[32]
port 102 nsew signal bidirectional
flabel metal2 s 16090 39200 16202 39800 0 FreeSans 448 90 0 0 io_out[33]
port 103 nsew signal bidirectional
flabel metal2 s 21886 39200 21998 39800 0 FreeSans 448 90 0 0 io_out[34]
port 104 nsew signal bidirectional
flabel metal2 s 38630 200 38742 800 0 FreeSans 448 90 0 0 io_out[35]
port 105 nsew signal bidirectional
flabel metal3 s 200 8788 800 9028 0 FreeSans 960 0 0 0 io_out[36]
port 106 nsew signal bidirectional
flabel metal3 s 39200 2668 39800 2908 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal bidirectional
flabel metal2 s 5786 200 5898 800 0 FreeSans 448 90 0 0 io_out[3]
port 108 nsew signal bidirectional
flabel metal3 s 200 21708 800 21948 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal bidirectional
flabel metal2 s 20598 39200 20710 39800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal bidirectional
flabel metal3 s 39200 17628 39800 17868 0 FreeSans 960 0 0 0 io_out[6]
port 111 nsew signal bidirectional
flabel metal3 s 39200 7428 39800 7668 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal bidirectional
flabel metal3 s 200 38028 800 38268 0 FreeSans 960 0 0 0 io_out[8]
port 113 nsew signal bidirectional
flabel metal3 s 39200 33268 39800 33508 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 115 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 115 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 116 nsew ground bidirectional
flabel metal2 s 12870 39200 12982 39800 0 FreeSans 448 90 0 0 wb_clk_i
port 117 nsew signal input
flabel metal3 s 39200 38708 39800 38948 0 FreeSans 960 0 0 0 wb_rst_i
port 118 nsew signal input
flabel metal3 s 200 28508 800 28748 0 FreeSans 960 0 0 0 wbs_ack_o
port 119 nsew signal bidirectional
flabel metal3 s 39200 25788 39800 26028 0 FreeSans 960 0 0 0 wbs_adr_i[0]
port 120 nsew signal input
flabel metal3 s 39200 32588 39800 32828 0 FreeSans 960 0 0 0 wbs_adr_i[10]
port 121 nsew signal input
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 wbs_adr_i[11]
port 122 nsew signal input
flabel metal2 s 1922 200 2034 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 123 nsew signal input
flabel metal2 s 15446 200 15558 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 124 nsew signal input
flabel metal3 s 39200 9468 39800 9708 0 FreeSans 960 0 0 0 wbs_adr_i[14]
port 125 nsew signal input
flabel metal2 s 19954 39200 20066 39800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 126 nsew signal input
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 127 nsew signal input
flabel metal3 s 39200 6748 39800 6988 0 FreeSans 960 0 0 0 wbs_adr_i[17]
port 128 nsew signal input
flabel metal2 s 37986 200 38098 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 129 nsew signal input
flabel metal3 s 200 35308 800 35548 0 FreeSans 960 0 0 0 wbs_adr_i[19]
port 130 nsew signal input
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 wbs_adr_i[1]
port 131 nsew signal input
flabel metal3 s 39200 21708 39800 21948 0 FreeSans 960 0 0 0 wbs_adr_i[20]
port 132 nsew signal input
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 wbs_adr_i[21]
port 133 nsew signal input
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 wbs_adr_i[22]
port 134 nsew signal input
flabel metal2 s 36054 200 36166 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 135 nsew signal input
flabel metal2 s 11582 39200 11694 39800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 136 nsew signal input
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 137 nsew signal input
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 wbs_adr_i[26]
port 138 nsew signal input
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 wbs_adr_i[27]
port 139 nsew signal input
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 wbs_adr_i[28]
port 140 nsew signal input
flabel metal2 s 10938 39200 11050 39800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 141 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 142 nsew signal input
flabel metal2 s 4498 39200 4610 39800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 143 nsew signal input
flabel metal3 s 39200 3348 39800 3588 0 FreeSans 960 0 0 0 wbs_adr_i[31]
port 144 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 145 nsew signal input
flabel metal3 s 39200 31228 39800 31468 0 FreeSans 960 0 0 0 wbs_adr_i[4]
port 146 nsew signal input
flabel metal3 s 200 4028 800 4268 0 FreeSans 960 0 0 0 wbs_adr_i[5]
port 147 nsew signal input
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 148 nsew signal input
flabel metal2 s 8362 39200 8474 39800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 149 nsew signal input
flabel metal2 s 31546 200 31658 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 150 nsew signal input
flabel metal3 s 200 24428 800 24668 0 FreeSans 960 0 0 0 wbs_adr_i[9]
port 151 nsew signal input
flabel metal2 s 31546 39200 31658 39800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 152 nsew signal input
flabel metal2 s 634 39200 746 39800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 153 nsew signal input
flabel metal2 s 9006 39200 9118 39800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 154 nsew signal input
flabel metal2 s 15446 39200 15558 39800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 155 nsew signal input
flabel metal2 s 14158 39200 14270 39800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 156 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 157 nsew signal input
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 158 nsew signal input
flabel metal3 s 200 10828 800 11068 0 FreeSans 960 0 0 0 wbs_dat_i[15]
port 159 nsew signal input
flabel metal2 s 18666 200 18778 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 160 nsew signal input
flabel metal3 s 39200 38028 39800 38268 0 FreeSans 960 0 0 0 wbs_dat_i[17]
port 161 nsew signal input
flabel metal2 s 1922 39200 2034 39800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 162 nsew signal input
flabel metal2 s 19310 39200 19422 39800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 163 nsew signal input
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 164 nsew signal input
flabel metal3 s 39200 14228 39800 14468 0 FreeSans 960 0 0 0 wbs_dat_i[20]
port 165 nsew signal input
flabel metal3 s 39200 29868 39800 30108 0 FreeSans 960 0 0 0 wbs_dat_i[21]
port 166 nsew signal input
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 wbs_dat_i[22]
port 167 nsew signal input
flabel metal3 s 39200 21028 39800 21268 0 FreeSans 960 0 0 0 wbs_dat_i[23]
port 168 nsew signal input
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 wbs_dat_i[24]
port 169 nsew signal input
flabel metal3 s 200 6068 800 6308 0 FreeSans 960 0 0 0 wbs_dat_i[25]
port 170 nsew signal input
flabel metal3 s 39200 35308 39800 35548 0 FreeSans 960 0 0 0 wbs_dat_i[26]
port 171 nsew signal input
flabel metal2 s 23174 39200 23286 39800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 172 nsew signal input
flabel metal2 s 10294 200 10406 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 173 nsew signal input
flabel metal3 s 39200 15588 39800 15828 0 FreeSans 960 0 0 0 wbs_dat_i[29]
port 174 nsew signal input
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 175 nsew signal input
flabel metal3 s 39200 5388 39800 5628 0 FreeSans 960 0 0 0 wbs_dat_i[30]
port 176 nsew signal input
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 wbs_dat_i[31]
port 177 nsew signal input
flabel metal2 s 35410 200 35522 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 178 nsew signal input
flabel metal2 s 5142 200 5254 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 179 nsew signal input
flabel metal2 s 16734 200 16846 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 180 nsew signal input
flabel metal3 s 39200 10148 39800 10388 0 FreeSans 960 0 0 0 wbs_dat_i[6]
port 181 nsew signal input
flabel metal3 s 39200 39388 39800 39628 0 FreeSans 960 0 0 0 wbs_dat_i[7]
port 182 nsew signal input
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 wbs_dat_i[8]
port 183 nsew signal input
flabel metal2 s 37342 200 37454 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 184 nsew signal input
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 wbs_dat_o[0]
port 185 nsew signal bidirectional
flabel metal3 s 39200 16268 39800 16508 0 FreeSans 960 0 0 0 wbs_dat_o[10]
port 186 nsew signal bidirectional
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 187 nsew signal bidirectional
flabel metal3 s 39200 30548 39800 30788 0 FreeSans 960 0 0 0 wbs_dat_o[12]
port 188 nsew signal bidirectional
flabel metal2 s 37342 39200 37454 39800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 189 nsew signal bidirectional
flabel metal3 s 39200 -52 39800 188 0 FreeSans 960 0 0 0 wbs_dat_o[14]
port 190 nsew signal bidirectional
flabel metal2 s 34766 39200 34878 39800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 191 nsew signal bidirectional
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 wbs_dat_o[16]
port 192 nsew signal bidirectional
flabel metal3 s 200 22388 800 22628 0 FreeSans 960 0 0 0 wbs_dat_o[17]
port 193 nsew signal bidirectional
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 194 nsew signal bidirectional
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 195 nsew signal bidirectional
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 196 nsew signal bidirectional
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 wbs_dat_o[20]
port 197 nsew signal bidirectional
flabel metal2 s 2566 39200 2678 39800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 198 nsew signal bidirectional
flabel metal2 s 17378 39200 17490 39800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 199 nsew signal bidirectional
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 wbs_dat_o[23]
port 200 nsew signal bidirectional
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 201 nsew signal bidirectional
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 202 nsew signal bidirectional
flabel metal2 s 25106 39200 25218 39800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 203 nsew signal bidirectional
flabel metal2 s 16734 39200 16846 39800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 204 nsew signal bidirectional
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 205 nsew signal bidirectional
flabel metal2 s 30902 39200 31014 39800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 206 nsew signal bidirectional
flabel metal3 s 39200 8108 39800 8348 0 FreeSans 960 0 0 0 wbs_dat_o[2]
port 207 nsew signal bidirectional
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 wbs_dat_o[30]
port 208 nsew signal bidirectional
flabel metal3 s 39200 28508 39800 28748 0 FreeSans 960 0 0 0 wbs_dat_o[31]
port 209 nsew signal bidirectional
flabel metal2 s 8362 200 8474 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 210 nsew signal bidirectional
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 211 nsew signal bidirectional
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 212 nsew signal bidirectional
flabel metal3 s 39200 27148 39800 27388 0 FreeSans 960 0 0 0 wbs_dat_o[6]
port 213 nsew signal bidirectional
flabel metal2 s 23174 200 23286 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 214 nsew signal bidirectional
flabel metal2 s 27682 39200 27794 39800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 215 nsew signal bidirectional
flabel metal2 s 27038 39200 27150 39800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 216 nsew signal bidirectional
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 wbs_sel_i[0]
port 217 nsew signal input
flabel metal2 s 5786 39200 5898 39800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 218 nsew signal input
flabel metal2 s 27038 200 27150 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 219 nsew signal input
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 wbs_sel_i[3]
port 220 nsew signal input
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 wbs_stb_i
port 221 nsew signal input
flabel metal3 s 39200 18308 39800 18548 0 FreeSans 960 0 0 0 wbs_we_i
port 222 nsew signal input
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel via1 20658 25942 20658 25942 0 _0000_
rlabel metal1 18216 27098 18216 27098 0 _0001_
rlabel metal2 12742 25670 12742 25670 0 _0002_
rlabel metal1 10610 29546 10610 29546 0 _0003_
rlabel metal1 10722 32402 10722 32402 0 _0004_
rlabel metal1 18818 23766 18818 23766 0 _0005_
rlabel metal1 15635 24106 15635 24106 0 _0006_
rlabel metal1 10518 24106 10518 24106 0 _0007_
rlabel metal1 10984 23086 10984 23086 0 _0008_
rlabel metal1 10150 20842 10150 20842 0 _0009_
rlabel metal2 12466 20706 12466 20706 0 _0010_
rlabel metal1 10978 17578 10978 17578 0 _0011_
rlabel metal1 10810 18394 10810 18394 0 _0012_
rlabel via1 11081 18734 11081 18734 0 _0013_
rlabel metal1 9798 22950 9798 22950 0 _0014_
rlabel metal1 14720 16762 14720 16762 0 _0015_
rlabel metal2 14674 34578 14674 34578 0 _0016_
rlabel metal2 14674 32674 14674 32674 0 _0017_
rlabel metal1 12599 32402 12599 32402 0 _0018_
rlabel metal1 13810 31790 13810 31790 0 _0019_
rlabel metal1 18533 29206 18533 29206 0 _0020_
rlabel metal1 21426 31790 21426 31790 0 _0021_
rlabel metal2 21298 33762 21298 33762 0 _0022_
rlabel metal1 21190 34986 21190 34986 0 _0023_
rlabel metal2 16974 35462 16974 35462 0 _0024_
rlabel via1 16601 32810 16601 32810 0 _0025_
rlabel metal1 21252 20026 21252 20026 0 _0026_
rlabel metal1 21742 28458 21742 28458 0 _0027_
rlabel metal1 24140 20910 24140 20910 0 _0028_
rlabel metal2 25530 33762 25530 33762 0 _0029_
rlabel metal1 21482 15980 21482 15980 0 _0030_
rlabel metal2 22494 24786 22494 24786 0 _0031_
rlabel metal1 23506 26350 23506 26350 0 _0032_
rlabel metal2 30130 31586 30130 31586 0 _0033_
rlabel metal1 29900 29818 29900 29818 0 _0034_
rlabel metal1 29067 25942 29067 25942 0 _0035_
rlabel metal2 28198 26384 28198 26384 0 _0036_
rlabel via1 24789 23698 24789 23698 0 _0037_
rlabel metal2 25530 27642 25530 27642 0 _0038_
rlabel metal2 29670 21794 29670 21794 0 _0039_
rlabel metal2 14582 18258 14582 18258 0 _0040_
rlabel metal2 17986 15844 17986 15844 0 _0041_
rlabel metal2 16238 14178 16238 14178 0 _0042_
rlabel metal1 20152 14382 20152 14382 0 _0043_
rlabel metal1 22820 13906 22820 13906 0 _0044_
rlabel metal1 15359 15470 15359 15470 0 _0045_
rlabel metal2 10258 14178 10258 14178 0 _0046_
rlabel via1 10713 13226 10713 13226 0 _0047_
rlabel metal1 14770 14314 14770 14314 0 _0048_
rlabel metal2 24426 21794 24426 21794 0 _0049_
rlabel via1 28009 21522 28009 21522 0 _0050_
rlabel metal1 27278 18156 27278 18156 0 _0051_
rlabel metal1 29435 19414 29435 19414 0 _0052_
rlabel metal1 27799 15402 27799 15402 0 _0053_
rlabel metal1 22627 22678 22627 22678 0 _0054_
rlabel metal1 25484 15130 25484 15130 0 _0055_
rlabel metal2 25162 13702 25162 13702 0 _0056_
rlabel metal2 2898 29801 2898 29801 0 _0057_
rlabel metal1 4830 37196 4830 37196 0 _0058_
rlabel metal1 37950 25874 37950 25874 0 _0059_
rlabel metal1 12098 3026 12098 3026 0 _0060_
rlabel metal1 37674 2448 37674 2448 0 _0061_
rlabel metal1 2346 4624 2346 4624 0 _0062_
rlabel metal1 4094 18258 4094 18258 0 _0063_
rlabel metal1 3266 2482 3266 2482 0 _0064_
rlabel metal1 2806 4556 2806 4556 0 _0065_
rlabel metal1 4784 6290 4784 6290 0 _0066_
rlabel metal1 2438 17680 2438 17680 0 _0067_
rlabel metal1 3956 24174 3956 24174 0 _0068_
rlabel metal1 37398 6290 37398 6290 0 _0069_
rlabel metal1 4554 16082 4554 16082 0 _0070_
rlabel metal1 24196 36006 24196 36006 0 _0071_
rlabel metal2 37490 4012 37490 4012 0 _0072_
rlabel metal1 37444 19822 37444 19822 0 _0073_
rlabel metal1 33856 23086 33856 23086 0 _0074_
rlabel metal2 2530 4352 2530 4352 0 _0075_
rlabel metal1 5198 3502 5198 3502 0 _0076_
rlabel metal1 25990 4046 25990 4046 0 _0077_
rlabel metal2 20746 24310 20746 24310 0 _0078_
rlabel metal2 18446 24990 18446 24990 0 _0079_
rlabel metal2 20838 29070 20838 29070 0 _0080_
rlabel metal1 19642 35088 19642 35088 0 _0081_
rlabel metal1 18814 31654 18814 31654 0 _0082_
rlabel via1 20102 33492 20102 33492 0 _0083_
rlabel metal2 29026 32606 29026 32606 0 _0084_
rlabel metal2 19642 32096 19642 32096 0 _0085_
rlabel metal1 18630 32198 18630 32198 0 _0086_
rlabel metal1 19826 32334 19826 32334 0 _0087_
rlabel metal1 20792 31790 20792 31790 0 _0088_
rlabel metal2 9982 31994 9982 31994 0 _0089_
rlabel metal1 8970 22678 8970 22678 0 _0090_
rlabel metal1 9200 23698 9200 23698 0 _0091_
rlabel metal1 11914 26928 11914 26928 0 _0092_
rlabel metal1 16100 20230 16100 20230 0 _0093_
rlabel metal1 17250 20434 17250 20434 0 _0094_
rlabel metal1 16928 24038 16928 24038 0 _0095_
rlabel metal1 13984 23562 13984 23562 0 _0096_
rlabel metal1 8464 29138 8464 29138 0 _0097_
rlabel metal2 19458 18462 19458 18462 0 _0098_
rlabel metal2 18722 17680 18722 17680 0 _0099_
rlabel metal1 18262 19686 18262 19686 0 _0100_
rlabel metal1 18262 20026 18262 20026 0 _0101_
rlabel metal2 14122 24004 14122 24004 0 _0102_
rlabel metal1 20424 31790 20424 31790 0 _0103_
rlabel metal1 20976 31858 20976 31858 0 _0104_
rlabel metal2 20102 21522 20102 21522 0 _0105_
rlabel metal1 12328 21318 12328 21318 0 _0106_
rlabel metal1 15456 21998 15456 21998 0 _0107_
rlabel metal1 20424 21522 20424 21522 0 _0108_
rlabel metal1 20102 28050 20102 28050 0 _0109_
rlabel metal1 20102 28118 20102 28118 0 _0110_
rlabel metal1 20148 27438 20148 27438 0 _0111_
rlabel metal1 35098 28084 35098 28084 0 _0112_
rlabel metal1 19412 32810 19412 32810 0 _0113_
rlabel metal2 19458 28492 19458 28492 0 _0114_
rlabel metal1 15594 21454 15594 21454 0 _0115_
rlabel metal2 14766 22508 14766 22508 0 _0116_
rlabel metal2 18262 23103 18262 23103 0 _0117_
rlabel metal1 17618 23562 17618 23562 0 _0118_
rlabel metal1 22678 31790 22678 31790 0 _0119_
rlabel metal2 19826 30056 19826 30056 0 _0120_
rlabel metal1 19918 27914 19918 27914 0 _0121_
rlabel metal1 15088 32402 15088 32402 0 _0122_
rlabel metal1 20010 27982 20010 27982 0 _0123_
rlabel metal2 19642 27642 19642 27642 0 _0124_
rlabel metal1 17825 28050 17825 28050 0 _0125_
rlabel metal1 27738 12716 27738 12716 0 _0126_
rlabel metal1 27508 21998 27508 21998 0 _0127_
rlabel metal2 24518 19516 24518 19516 0 _0128_
rlabel metal2 25990 17850 25990 17850 0 _0129_
rlabel metal1 30314 16014 30314 16014 0 _0130_
rlabel metal1 26818 17306 26818 17306 0 _0131_
rlabel metal1 26956 33014 26956 33014 0 _0132_
rlabel metal2 25898 31042 25898 31042 0 _0133_
rlabel metal1 28014 30158 28014 30158 0 _0134_
rlabel metal1 29532 30906 29532 30906 0 _0135_
rlabel metal2 28566 28050 28566 28050 0 _0136_
rlabel metal1 27692 27574 27692 27574 0 _0137_
rlabel metal1 26818 27302 26818 27302 0 _0138_
rlabel metal2 23138 17374 23138 17374 0 _0139_
rlabel metal2 13478 19040 13478 19040 0 _0140_
rlabel metal1 15916 26010 15916 26010 0 _0141_
rlabel metal1 15548 25466 15548 25466 0 _0142_
rlabel metal1 15732 25806 15732 25806 0 _0143_
rlabel metal2 10810 26452 10810 26452 0 _0144_
rlabel metal1 12098 28730 12098 28730 0 _0145_
rlabel metal1 14168 29478 14168 29478 0 _0146_
rlabel metal1 14444 29070 14444 29070 0 _0147_
rlabel metal1 14306 30022 14306 30022 0 _0148_
rlabel metal2 13294 28764 13294 28764 0 _0149_
rlabel metal2 13386 27778 13386 27778 0 _0150_
rlabel metal1 10994 27506 10994 27506 0 _0151_
rlabel metal2 11178 27812 11178 27812 0 _0152_
rlabel metal1 12374 25976 12374 25976 0 _0153_
rlabel metal2 14306 30260 14306 30260 0 _0154_
rlabel metal1 8786 30260 8786 30260 0 _0155_
rlabel metal2 9706 31756 9706 31756 0 _0156_
rlabel metal2 9062 30328 9062 30328 0 _0157_
rlabel metal1 9200 30158 9200 30158 0 _0158_
rlabel metal1 9476 27438 9476 27438 0 _0159_
rlabel metal2 10902 26554 10902 26554 0 _0160_
rlabel metal1 11454 26010 11454 26010 0 _0161_
rlabel metal1 9660 26350 9660 26350 0 _0162_
rlabel metal1 8924 26554 8924 26554 0 _0163_
rlabel metal1 9384 25874 9384 25874 0 _0164_
rlabel metal2 9430 26588 9430 26588 0 _0165_
rlabel metal2 9614 27030 9614 27030 0 _0166_
rlabel metal1 10442 27574 10442 27574 0 _0167_
rlabel metal1 12282 28152 12282 28152 0 _0168_
rlabel metal1 16859 18258 16859 18258 0 _0169_
rlabel metal1 15088 32198 15088 32198 0 _0170_
rlabel metal2 15778 28220 15778 28220 0 _0171_
rlabel metal2 15594 28492 15594 28492 0 _0172_
rlabel metal1 9246 25942 9246 25942 0 _0173_
rlabel metal1 8740 26010 8740 26010 0 _0174_
rlabel metal1 8510 29614 8510 29614 0 _0175_
rlabel metal1 8694 28526 8694 28526 0 _0176_
rlabel metal2 7866 28764 7866 28764 0 _0177_
rlabel metal2 8786 28186 8786 28186 0 _0178_
rlabel metal1 15042 28050 15042 28050 0 _0179_
rlabel metal1 17250 28152 17250 28152 0 _0180_
rlabel metal1 17066 27880 17066 27880 0 _0181_
rlabel metal2 15502 28220 15502 28220 0 _0182_
rlabel metal1 16100 27642 16100 27642 0 _0183_
rlabel metal1 5589 26962 5589 26962 0 _0184_
rlabel metal1 17296 32198 17296 32198 0 _0185_
rlabel metal1 16146 31790 16146 31790 0 _0186_
rlabel via1 17894 22073 17894 22073 0 _0187_
rlabel metal1 21068 19278 21068 19278 0 _0188_
rlabel metal2 15134 21692 15134 21692 0 _0189_
rlabel metal1 17526 21556 17526 21556 0 _0190_
rlabel metal1 17756 17238 17756 17238 0 _0191_
rlabel metal1 18400 31790 18400 31790 0 _0192_
rlabel metal1 17894 19210 17894 19210 0 _0193_
rlabel metal2 17434 21590 17434 21590 0 _0194_
rlabel metal1 16606 22406 16606 22406 0 _0195_
rlabel metal2 13294 20876 13294 20876 0 _0196_
rlabel metal1 15226 20570 15226 20570 0 _0197_
rlabel metal2 17802 24174 17802 24174 0 _0198_
rlabel metal1 18170 25976 18170 25976 0 _0199_
rlabel metal1 18032 16150 18032 16150 0 _0200_
rlabel metal2 11914 28764 11914 28764 0 _0201_
rlabel metal1 19550 19414 19550 19414 0 _0202_
rlabel metal1 19872 25466 19872 25466 0 _0203_
rlabel metal2 12374 26860 12374 26860 0 _0204_
rlabel metal2 17434 26792 17434 26792 0 _0205_
rlabel metal1 17848 26962 17848 26962 0 _0206_
rlabel metal2 12834 26758 12834 26758 0 _0207_
rlabel metal1 12450 26282 12450 26282 0 _0208_
rlabel metal2 12926 25738 12926 25738 0 _0209_
rlabel metal2 11822 30294 11822 30294 0 _0210_
rlabel metal2 11914 29648 11914 29648 0 _0211_
rlabel metal1 10902 29274 10902 29274 0 _0212_
rlabel metal2 10442 32436 10442 32436 0 _0213_
rlabel metal1 17710 24208 17710 24208 0 _0214_
rlabel metal1 17618 24684 17618 24684 0 _0215_
rlabel metal1 10258 23052 10258 23052 0 _0216_
rlabel metal2 16698 24616 16698 24616 0 _0217_
rlabel metal1 9338 24378 9338 24378 0 _0218_
rlabel metal1 20286 34170 20286 34170 0 _0219_
rlabel metal1 9936 24582 9936 24582 0 _0220_
rlabel via1 9798 23698 9798 23698 0 _0221_
rlabel metal1 10028 24786 10028 24786 0 _0222_
rlabel metal1 9522 23494 9522 23494 0 _0223_
rlabel metal2 9062 23868 9062 23868 0 _0224_
rlabel metal2 9154 21318 9154 21318 0 _0225_
rlabel metal1 16146 19210 16146 19210 0 _0226_
rlabel metal1 9706 21556 9706 21556 0 _0227_
rlabel metal1 9798 20400 9798 20400 0 _0228_
rlabel metal1 9108 20434 9108 20434 0 _0229_
rlabel metal1 9430 18054 9430 18054 0 _0230_
rlabel metal1 10028 17646 10028 17646 0 _0231_
rlabel metal2 10350 19108 10350 19108 0 _0232_
rlabel metal1 10534 18292 10534 18292 0 _0233_
rlabel metal1 9476 22474 9476 22474 0 _0234_
rlabel metal1 14950 16558 14950 16558 0 _0235_
rlabel metal1 9476 22542 9476 22542 0 _0236_
rlabel metal2 10534 16320 10534 16320 0 _0237_
rlabel metal2 11822 16252 11822 16252 0 _0238_
rlabel metal2 10350 14246 10350 14246 0 _0239_
rlabel metal1 13156 14790 13156 14790 0 _0240_
rlabel metal2 13018 17612 13018 17612 0 _0241_
rlabel metal2 9154 14722 9154 14722 0 _0242_
rlabel metal1 12790 16558 12790 16558 0 _0243_
rlabel metal1 10672 16490 10672 16490 0 _0244_
rlabel metal2 12926 16898 12926 16898 0 _0245_
rlabel metal1 16698 18598 16698 18598 0 _0246_
rlabel metal1 17020 18326 17020 18326 0 _0247_
rlabel metal1 17378 18224 17378 18224 0 _0248_
rlabel via1 20026 14994 20026 14994 0 _0249_
rlabel metal2 18170 18088 18170 18088 0 _0250_
rlabel metal1 17296 18394 17296 18394 0 _0251_
rlabel metal2 20194 14144 20194 14144 0 _0252_
rlabel metal1 17572 16762 17572 16762 0 _0253_
rlabel metal1 20010 11628 20010 11628 0 _0254_
rlabel metal2 17342 19516 17342 19516 0 _0255_
rlabel metal2 16330 18496 16330 18496 0 _0256_
rlabel metal1 17526 18938 17526 18938 0 _0257_
rlabel metal2 18354 19618 18354 19618 0 _0258_
rlabel metal1 22402 11764 22402 11764 0 _0259_
rlabel metal1 16833 19812 16833 19812 0 _0260_
rlabel metal2 17158 19584 17158 19584 0 _0261_
rlabel metal2 13570 16898 13570 16898 0 _0262_
rlabel metal2 12466 15164 12466 15164 0 _0263_
rlabel metal1 13156 15130 13156 15130 0 _0264_
rlabel metal1 13340 16762 13340 16762 0 _0265_
rlabel metal1 14260 16626 14260 16626 0 _0266_
rlabel metal1 11362 16558 11362 16558 0 _0267_
rlabel metal1 14398 16524 14398 16524 0 _0268_
rlabel metal1 19964 34510 19964 34510 0 _0269_
rlabel metal2 14490 34170 14490 34170 0 _0270_
rlabel metal2 14858 32844 14858 32844 0 _0271_
rlabel metal2 15226 30498 15226 30498 0 _0272_
rlabel metal1 15272 31382 15272 31382 0 _0273_
rlabel metal1 13570 32878 13570 32878 0 _0274_
rlabel metal2 20654 30328 20654 30328 0 _0275_
rlabel metal1 18814 30668 18814 30668 0 _0276_
rlabel metal2 18170 31586 18170 31586 0 _0277_
rlabel metal1 19182 35122 19182 35122 0 _0278_
rlabel metal2 21022 33490 21022 33490 0 _0279_
rlabel metal2 21114 33660 21114 33660 0 _0280_
rlabel metal1 20424 34578 20424 34578 0 _0281_
rlabel metal2 21022 34884 21022 34884 0 _0282_
rlabel metal2 18170 34748 18170 34748 0 _0283_
rlabel metal2 18446 34408 18446 34408 0 _0284_
rlabel metal2 17618 34884 17618 34884 0 _0285_
rlabel metal1 17020 33626 17020 33626 0 _0286_
rlabel metal1 22724 18870 22724 18870 0 _0287_
rlabel metal2 24058 20094 24058 20094 0 _0288_
rlabel metal2 23230 19788 23230 19788 0 _0289_
rlabel metal1 24334 17204 24334 17204 0 _0290_
rlabel metal1 23966 18598 23966 18598 0 _0291_
rlabel metal2 20838 19108 20838 19108 0 _0292_
rlabel metal1 19366 20502 19366 20502 0 _0293_
rlabel metal2 19366 20876 19366 20876 0 _0294_
rlabel metal2 18538 21420 18538 21420 0 _0295_
rlabel metal1 18584 20502 18584 20502 0 _0296_
rlabel metal2 18998 20604 18998 20604 0 _0297_
rlabel metal1 20654 19822 20654 19822 0 _0298_
rlabel metal1 20654 19992 20654 19992 0 _0299_
rlabel metal2 20010 18666 20010 18666 0 _0300_
rlabel metal2 20746 19516 20746 19516 0 _0301_
rlabel metal1 19918 19176 19918 19176 0 _0302_
rlabel metal1 25162 17102 25162 17102 0 _0303_
rlabel metal2 21206 17442 21206 17442 0 _0304_
rlabel metal1 20792 18054 20792 18054 0 _0305_
rlabel metal2 20654 18564 20654 18564 0 _0306_
rlabel metal2 23598 18870 23598 18870 0 _0307_
rlabel metal1 22724 19142 22724 19142 0 _0308_
rlabel metal1 23460 19346 23460 19346 0 _0309_
rlabel metal2 23506 18700 23506 18700 0 _0310_
rlabel metal1 23828 17306 23828 17306 0 _0311_
rlabel metal1 23000 18394 23000 18394 0 _0312_
rlabel metal2 20378 18258 20378 18258 0 _0313_
rlabel metal2 20194 19176 20194 19176 0 _0314_
rlabel metal1 20792 19482 20792 19482 0 _0315_
rlabel metal1 21114 28458 21114 28458 0 _0316_
rlabel metal2 21206 28730 21206 28730 0 _0317_
rlabel metal1 21804 16558 21804 16558 0 _0318_
rlabel metal1 20378 22202 20378 22202 0 _0319_
rlabel metal2 27646 19278 27646 19278 0 _0320_
rlabel metal1 21643 21522 21643 21522 0 _0321_
rlabel metal1 20930 22542 20930 22542 0 _0322_
rlabel metal1 23368 30226 23368 30226 0 _0323_
rlabel metal2 23138 30430 23138 30430 0 _0324_
rlabel metal2 22126 30260 22126 30260 0 _0325_
rlabel metal2 22402 30362 22402 30362 0 _0326_
rlabel metal1 24978 32266 24978 32266 0 _0327_
rlabel metal2 27278 33796 27278 33796 0 _0328_
rlabel metal1 28014 33932 28014 33932 0 _0329_
rlabel metal2 27186 33116 27186 33116 0 _0330_
rlabel metal1 27968 31450 27968 31450 0 _0331_
rlabel metal1 27968 31994 27968 31994 0 _0332_
rlabel metal1 27324 32878 27324 32878 0 _0333_
rlabel metal2 25254 32130 25254 32130 0 _0334_
rlabel metal1 24610 31688 24610 31688 0 _0335_
rlabel metal1 24840 31994 24840 31994 0 _0336_
rlabel metal1 24518 30090 24518 30090 0 _0337_
rlabel metal1 25162 31994 25162 31994 0 _0338_
rlabel metal1 24610 32538 24610 32538 0 _0339_
rlabel metal1 25760 25262 25760 25262 0 _0340_
rlabel metal1 24656 33286 24656 33286 0 _0341_
rlabel metal2 27462 32929 27462 32929 0 _0342_
rlabel metal1 26220 32878 26220 32878 0 _0343_
rlabel metal1 26496 33082 26496 33082 0 _0344_
rlabel metal1 27784 31790 27784 31790 0 _0345_
rlabel metal1 28566 31824 28566 31824 0 _0346_
rlabel metal2 27094 32164 27094 32164 0 _0347_
rlabel metal2 28198 33116 28198 33116 0 _0348_
rlabel metal2 27554 32572 27554 32572 0 _0349_
rlabel metal2 26082 32708 26082 32708 0 _0350_
rlabel metal1 25530 32980 25530 32980 0 _0351_
rlabel metal1 24794 31450 24794 31450 0 _0352_
rlabel metal2 25622 31110 25622 31110 0 _0353_
rlabel metal2 25162 32130 25162 32130 0 _0354_
rlabel metal1 25714 32776 25714 32776 0 _0355_
rlabel metal2 25622 33286 25622 33286 0 _0356_
rlabel metal1 25116 33490 25116 33490 0 _0357_
rlabel metal1 15640 13906 15640 13906 0 _0358_
rlabel metal1 21344 16762 21344 16762 0 _0359_
rlabel metal2 21298 16252 21298 16252 0 _0360_
rlabel metal1 15364 21658 15364 21658 0 _0361_
rlabel metal1 16698 21862 16698 21862 0 _0362_
rlabel metal2 17802 15079 17802 15079 0 _0363_
rlabel metal1 23736 21998 23736 21998 0 _0364_
rlabel viali 22959 24174 22959 24174 0 _0365_
rlabel metal2 29854 14110 29854 14110 0 _0366_
rlabel metal1 27646 17714 27646 17714 0 _0367_
rlabel metal2 24702 26554 24702 26554 0 _0368_
rlabel metal1 20286 23188 20286 23188 0 _0369_
rlabel metal2 27186 21794 27186 21794 0 _0370_
rlabel metal2 23046 27642 23046 27642 0 _0371_
rlabel metal2 24058 27642 24058 27642 0 _0372_
rlabel via1 22957 27302 22957 27302 0 _0373_
rlabel metal2 23506 27404 23506 27404 0 _0374_
rlabel metal1 24472 26350 24472 26350 0 _0375_
rlabel metal1 24932 13294 24932 13294 0 _0376_
rlabel metal2 31786 27540 31786 27540 0 _0377_
rlabel metal1 32016 27438 32016 27438 0 _0378_
rlabel metal2 32338 28866 32338 28866 0 _0379_
rlabel metal2 32522 28526 32522 28526 0 _0380_
rlabel metal1 31694 29614 31694 29614 0 _0381_
rlabel via1 30774 20230 30774 20230 0 _0382_
rlabel metal2 30590 30566 30590 30566 0 _0383_
rlabel metal2 30406 28220 30406 28220 0 _0384_
rlabel metal1 31418 28662 31418 28662 0 _0385_
rlabel metal1 31096 29206 31096 29206 0 _0386_
rlabel metal2 31050 28594 31050 28594 0 _0387_
rlabel metal2 32706 29750 32706 29750 0 _0388_
rlabel metal1 32614 30124 32614 30124 0 _0389_
rlabel metal1 31050 30090 31050 30090 0 _0390_
rlabel metal2 29946 29818 29946 29818 0 _0391_
rlabel metal1 30544 15334 30544 15334 0 _0392_
rlabel metal1 30958 28084 30958 28084 0 _0393_
rlabel metal2 31510 26554 31510 26554 0 _0394_
rlabel metal1 31372 25262 31372 25262 0 _0395_
rlabel metal1 30590 24786 30590 24786 0 _0396_
rlabel metal1 30682 24582 30682 24582 0 _0397_
rlabel metal1 29440 24650 29440 24650 0 _0398_
rlabel metal2 29118 25024 29118 25024 0 _0399_
rlabel metal2 29762 24582 29762 24582 0 _0400_
rlabel metal2 28658 24412 28658 24412 0 _0401_
rlabel metal2 29210 24004 29210 24004 0 _0402_
rlabel metal1 28152 24242 28152 24242 0 _0403_
rlabel metal2 28934 24582 28934 24582 0 _0404_
rlabel metal2 25162 24412 25162 24412 0 _0405_
rlabel metal1 27554 25262 27554 25262 0 _0406_
rlabel metal1 26864 24582 26864 24582 0 _0407_
rlabel metal1 26588 24718 26588 24718 0 _0408_
rlabel metal1 25622 25840 25622 25840 0 _0409_
rlabel metal2 26542 24582 26542 24582 0 _0410_
rlabel metal1 25300 24378 25300 24378 0 _0411_
rlabel metal2 25714 27200 25714 27200 0 _0412_
rlabel metal2 26358 26384 26358 26384 0 _0413_
rlabel metal1 26082 25942 26082 25942 0 _0414_
rlabel metal1 26404 26554 26404 26554 0 _0415_
rlabel metal1 26036 25670 26036 25670 0 _0416_
rlabel metal2 25806 26758 25806 26758 0 _0417_
rlabel metal1 16790 14994 16790 14994 0 _0418_
rlabel metal1 26956 25330 26956 25330 0 _0419_
rlabel metal2 27094 25738 27094 25738 0 _0420_
rlabel metal2 31878 24242 31878 24242 0 _0421_
rlabel metal1 31786 23188 31786 23188 0 _0422_
rlabel metal2 31050 22780 31050 22780 0 _0423_
rlabel metal1 30084 21522 30084 21522 0 _0424_
rlabel metal1 15916 12682 15916 12682 0 _0425_
rlabel metal1 12282 2618 12282 2618 0 _0426_
rlabel metal1 17434 12308 17434 12308 0 _0427_
rlabel metal1 17572 13294 17572 13294 0 _0428_
rlabel metal2 17342 17476 17342 17476 0 _0429_
rlabel metal2 21850 11730 21850 11730 0 _0430_
rlabel metal1 17618 15436 17618 15436 0 _0431_
rlabel metal1 17526 15504 17526 15504 0 _0432_
rlabel metal2 16146 13328 16146 13328 0 _0433_
rlabel metal1 18354 12206 18354 12206 0 _0434_
rlabel metal1 13478 11594 13478 11594 0 _0435_
rlabel metal2 19826 11458 19826 11458 0 _0436_
rlabel metal1 18492 12342 18492 12342 0 _0437_
rlabel metal1 18354 12410 18354 12410 0 _0438_
rlabel metal2 17986 13158 17986 13158 0 _0439_
rlabel metal2 16974 13702 16974 13702 0 _0440_
rlabel metal1 20286 12852 20286 12852 0 _0441_
rlabel metal1 19826 12818 19826 12818 0 _0442_
rlabel metal2 20010 12512 20010 12512 0 _0443_
rlabel metal1 22218 11594 22218 11594 0 _0444_
rlabel metal1 20194 12240 20194 12240 0 _0445_
rlabel metal1 20516 12410 20516 12410 0 _0446_
rlabel metal1 19688 14994 19688 14994 0 _0447_
rlabel metal1 22540 13498 22540 13498 0 _0448_
rlabel via1 21206 11526 21206 11526 0 _0449_
rlabel metal1 21988 11866 21988 11866 0 _0450_
rlabel metal2 21482 11900 21482 11900 0 _0451_
rlabel metal2 22126 13396 22126 13396 0 _0452_
rlabel metal1 18860 14246 18860 14246 0 _0453_
rlabel metal1 15962 12614 15962 12614 0 _0454_
rlabel metal1 16744 12206 16744 12206 0 _0455_
rlabel metal1 16146 11730 16146 11730 0 _0456_
rlabel metal1 15962 11696 15962 11696 0 _0457_
rlabel metal1 16238 11866 16238 11866 0 _0458_
rlabel metal1 17296 16082 17296 16082 0 _0459_
rlabel metal2 16882 16422 16882 16422 0 _0460_
rlabel metal2 15686 16252 15686 16252 0 _0461_
rlabel metal1 13984 11662 13984 11662 0 _0462_
rlabel metal2 12742 11322 12742 11322 0 _0463_
rlabel metal2 11270 13022 11270 13022 0 _0464_
rlabel metal2 9522 13090 9522 13090 0 _0465_
rlabel metal1 10028 13498 10028 13498 0 _0466_
rlabel metal2 11822 11900 11822 11900 0 _0467_
rlabel metal1 10626 12240 10626 12240 0 _0468_
rlabel metal1 10580 12410 10580 12410 0 _0469_
rlabel metal1 14996 13974 14996 13974 0 _0470_
rlabel metal1 12788 12206 12788 12206 0 _0471_
rlabel metal1 13202 12410 13202 12410 0 _0472_
rlabel metal1 14076 13498 14076 13498 0 _0473_
rlabel metal2 14214 14518 14214 14518 0 _0474_
rlabel metal2 23966 21692 23966 21692 0 _0475_
rlabel metal1 28152 20774 28152 20774 0 _0476_
rlabel metal1 27370 20264 27370 20264 0 _0477_
rlabel metal1 27822 20570 27822 20570 0 _0478_
rlabel metal1 27600 20026 27600 20026 0 _0479_
rlabel metal2 27002 20026 27002 20026 0 _0480_
rlabel metal1 27554 19958 27554 19958 0 _0481_
rlabel metal1 27508 17850 27508 17850 0 _0482_
rlabel metal1 28566 18802 28566 18802 0 _0483_
rlabel metal1 31878 18768 31878 18768 0 _0484_
rlabel via1 32062 18258 32062 18258 0 _0485_
rlabel metal1 28520 17646 28520 17646 0 _0486_
rlabel metal2 28290 18122 28290 18122 0 _0487_
rlabel metal1 27968 17850 27968 17850 0 _0488_
rlabel metal2 31142 20230 31142 20230 0 _0489_
rlabel metal1 31234 20298 31234 20298 0 _0490_
rlabel metal2 31694 18564 31694 18564 0 _0491_
rlabel metal2 31878 19414 31878 19414 0 _0492_
rlabel metal2 31694 20196 31694 20196 0 _0493_
rlabel metal2 29946 20026 29946 20026 0 _0494_
rlabel metal1 31096 17714 31096 17714 0 _0495_
rlabel metal2 30314 17408 30314 17408 0 _0496_
rlabel metal1 31326 16048 31326 16048 0 _0497_
rlabel metal1 30176 16422 30176 16422 0 _0498_
rlabel metal2 30222 15402 30222 15402 0 _0499_
rlabel metal2 30682 15300 30682 15300 0 _0500_
rlabel metal1 29624 15470 29624 15470 0 _0501_
rlabel via1 28290 15946 28290 15946 0 _0502_
rlabel metal1 30820 16762 30820 16762 0 _0503_
rlabel metal2 28382 16796 28382 16796 0 _0504_
rlabel metal2 27922 17833 27922 17833 0 _0505_
rlabel metal1 25944 21998 25944 21998 0 _0506_
rlabel metal1 22448 23086 22448 23086 0 _0507_
rlabel metal1 27876 12206 27876 12206 0 _0508_
rlabel metal1 28198 12614 28198 12614 0 _0509_
rlabel metal1 28060 12410 28060 12410 0 _0510_
rlabel metal1 28750 16082 28750 16082 0 _0511_
rlabel metal1 28566 13838 28566 13838 0 _0512_
rlabel metal2 27922 14212 27922 14212 0 _0513_
rlabel metal2 27278 14790 27278 14790 0 _0514_
rlabel metal1 26910 12818 26910 12818 0 _0515_
rlabel metal1 25530 12716 25530 12716 0 _0516_
rlabel metal1 26680 12954 26680 12954 0 _0517_
rlabel metal1 25668 13294 25668 13294 0 _0518_
rlabel metal2 2806 28900 2806 28900 0 _0519_
rlabel metal2 2254 14484 2254 14484 0 _0520_
rlabel metal2 28106 3230 28106 3230 0 _0521_
rlabel metal2 37582 7650 37582 7650 0 _0522_
rlabel metal1 8464 2618 8464 2618 0 _0523_
rlabel metal1 12742 2958 12742 2958 0 _0524_
rlabel metal1 22172 2618 22172 2618 0 _0525_
rlabel metal2 37582 27234 37582 27234 0 _0526_
rlabel metal1 23782 2618 23782 2618 0 _0527_
rlabel metal2 28014 35428 28014 35428 0 _0528_
rlabel metal1 26864 36074 26864 36074 0 _0529_
rlabel metal2 36662 15708 36662 15708 0 _0530_
rlabel metal2 9062 3230 9062 3230 0 _0531_
rlabel metal1 37904 30362 37904 30362 0 _0532_
rlabel metal1 37398 36074 37398 36074 0 _0533_
rlabel metal1 37214 2346 37214 2346 0 _0534_
rlabel metal1 34914 35258 34914 35258 0 _0535_
rlabel metal2 3266 21148 3266 21148 0 _0536_
rlabel metal2 3542 22814 3542 22814 0 _0537_
rlabel metal2 5750 4012 5750 4012 0 _0538_
rlabel metal2 2254 4964 2254 4964 0 _0539_
rlabel metal1 2116 27642 2116 27642 0 _0540_
rlabel metal1 3634 31450 3634 31450 0 _0541_
rlabel metal2 18722 36652 18722 36652 0 _0542_
rlabel metal2 2714 20196 2714 20196 0 _0543_
rlabel metal2 7498 2788 7498 2788 0 _0544_
rlabel metal1 3772 2346 3772 2346 0 _0545_
rlabel metal1 24242 35802 24242 35802 0 _0546_
rlabel metal2 14674 36958 14674 36958 0 _0547_
rlabel metal1 19872 3094 19872 3094 0 _0548_
rlabel metal1 31464 35802 31464 35802 0 _0549_
rlabel metal2 1794 31212 1794 31212 0 _0550_
rlabel metal1 38180 28730 38180 28730 0 _0551_
rlabel metal1 3312 35802 3312 35802 0 _0552_
rlabel metal2 3818 4318 3818 4318 0 _0553_
rlabel metal2 38134 12444 38134 12444 0 _0554_
rlabel metal2 5566 6562 5566 6562 0 _0555_
rlabel metal2 2438 21794 2438 21794 0 _0556_
rlabel metal2 19918 36516 19918 36516 0 _0557_
rlabel metal2 37582 17442 37582 17442 0 _0558_
rlabel metal1 38180 7174 38180 7174 0 _0559_
rlabel metal1 2116 35802 2116 35802 0 _0560_
rlabel metal1 36616 32538 36616 32538 0 _0561_
rlabel metal2 3542 4318 3542 4318 0 _0562_
rlabel metal1 20884 2618 20884 2618 0 _0563_
rlabel metal1 2208 17850 2208 17850 0 _0564_
rlabel metal2 23782 34068 23782 34068 0 _0565_
rlabel metal2 36018 28322 36018 28322 0 _0566_
rlabel metal2 4094 25619 4094 25619 0 _0567_
rlabel metal2 4094 24548 4094 24548 0 _0568_
rlabel metal2 14398 24004 14398 24004 0 _0569_
rlabel metal1 23690 9486 23690 9486 0 _0570_
rlabel metal2 33810 33966 33810 33966 0 _0571_
rlabel metal2 3266 14994 3266 14994 0 _0572_
rlabel metal1 29670 3434 29670 3434 0 _0573_
rlabel metal1 35788 35258 35788 35258 0 _0574_
rlabel metal1 26726 35734 26726 35734 0 _0575_
rlabel metal2 38134 24412 38134 24412 0 _0576_
rlabel metal1 4554 29818 4554 29818 0 _0577_
rlabel metal2 38134 5916 38134 5916 0 _0578_
rlabel metal2 36662 16796 36662 16796 0 _0579_
rlabel metal1 24012 36346 24012 36346 0 _0580_
rlabel metal1 29164 35258 29164 35258 0 _0581_
rlabel metal1 3036 10778 3036 10778 0 _0582_
rlabel metal1 25806 35802 25806 35802 0 _0583_
rlabel metal2 9430 36516 9430 36516 0 _0584_
rlabel metal1 15042 35802 15042 35802 0 _0585_
rlabel metal1 21160 35802 21160 35802 0 _0586_
rlabel metal1 35742 3434 35742 3434 0 _0587_
rlabel metal2 3266 9180 3266 9180 0 _0588_
rlabel metal1 36754 4012 36754 4012 0 _0589_
rlabel metal2 26082 3740 26082 3740 0 _0590_
rlabel metal1 37812 3162 37812 3162 0 _0591_
rlabel metal2 3266 30362 3266 30362 0 _0592_
rlabel metal2 6486 36516 6486 36516 0 _0593_
rlabel metal2 38134 11356 38134 11356 0 _0594_
rlabel metal2 2070 33694 2070 33694 0 _0595_
rlabel metal1 3956 35802 3956 35802 0 _0596_
rlabel metal2 35374 34680 35374 34680 0 _0597_
rlabel metal2 38134 19244 38134 19244 0 _0598_
rlabel metal2 3542 17374 3542 17374 0 _0599_
rlabel metal1 29992 35802 29992 35802 0 _0600_
rlabel metal2 34178 3230 34178 3230 0 _0601_
rlabel metal2 30130 36210 30130 36210 0 _0602_
rlabel metal1 33994 23290 33994 23290 0 _0603_
rlabel metal2 34086 31518 34086 31518 0 _0604_
rlabel metal1 33442 21454 33442 21454 0 _0605_
rlabel metal2 11638 11356 11638 11356 0 _0606_
rlabel metal1 18584 10234 18584 10234 0 _0607_
rlabel metal2 32430 33762 32430 33762 0 _0608_
rlabel metal2 2438 6562 2438 6562 0 _0609_
rlabel metal1 2898 2618 2898 2618 0 _0610_
rlabel metal2 10626 3740 10626 3740 0 _0611_
rlabel metal2 36754 35054 36754 35054 0 _0612_
rlabel metal1 32154 36822 32154 36822 0 _0613_
rlabel metal2 4370 3230 4370 3230 0 _0614_
rlabel metal1 11546 2346 11546 2346 0 _0615_
rlabel metal2 38134 22236 38134 22236 0 _0616_
rlabel metal1 24840 2482 24840 2482 0 _0617_
rlabel metal2 1794 12444 1794 12444 0 _0618_
rlabel metal1 18906 35802 18906 35802 0 _0619_
rlabel metal2 4370 36958 4370 36958 0 _0620_
rlabel metal2 38226 37026 38226 37026 0 _0621_
rlabel metal2 22310 36958 22310 36958 0 _0622_
rlabel metal2 36846 33762 36846 33762 0 _0623_
rlabel metal2 37582 34850 37582 34850 0 _0624_
rlabel metal1 4600 28594 4600 28594 0 _0625_
rlabel metal1 32890 35258 32890 35258 0 _0626_
rlabel metal2 38134 25500 38134 25500 0 _0627_
rlabel metal1 874 37230 874 37230 0 active
rlabel metal2 4002 26588 4002 26588 0 adapter.blue
rlabel metal1 21206 21998 21206 21998 0 adapter.debug_design_reset
rlabel metal1 31556 28526 31556 28526 0 adapter.game.ballDirX
rlabel metal1 26312 19822 26312 19822 0 adapter.game.ballDirY
rlabel metal2 24058 25908 24058 25908 0 adapter.game.ballX\[0\]
rlabel metal2 22770 29104 22770 29104 0 adapter.game.ballX\[1\]
rlabel metal1 23598 31824 23598 31824 0 adapter.game.ballX\[2\]
rlabel metal1 28934 29546 28934 29546 0 adapter.game.ballX\[3\]
rlabel metal1 30130 25772 30130 25772 0 adapter.game.ballX\[4\]
rlabel metal1 28880 29478 28880 29478 0 adapter.game.ballX\[5\]
rlabel metal1 27370 33456 27370 33456 0 adapter.game.ballX\[6\]
rlabel metal2 26542 29886 26542 29886 0 adapter.game.ballX\[7\]
rlabel metal2 24794 26061 24794 26061 0 adapter.game.ballX\[8\]
rlabel metal1 26358 20978 26358 20978 0 adapter.game.ballY\[0\]
rlabel metal1 19412 21522 19412 21522 0 adapter.game.ballY\[1\]
rlabel metal1 31878 17816 31878 17816 0 adapter.game.ballY\[2\]
rlabel metal2 30130 19686 30130 19686 0 adapter.game.ballY\[3\]
rlabel metal1 25530 18802 25530 18802 0 adapter.game.ballY\[4\]
rlabel metal1 23184 21454 23184 21454 0 adapter.game.ballY\[5\]
rlabel metal2 23598 15572 23598 15572 0 adapter.game.ballY\[6\]
rlabel metal2 21022 17408 21022 17408 0 adapter.game.ballY\[7\]
rlabel metal2 35282 28356 35282 28356 0 adapter.game.green
rlabel metal1 15410 34034 15410 34034 0 adapter.game.h\[0\]
rlabel metal1 17204 31790 17204 31790 0 adapter.game.h\[1\]
rlabel metal1 13846 30226 13846 30226 0 adapter.game.h\[2\]
rlabel metal1 9844 31722 9844 31722 0 adapter.game.h\[3\]
rlabel metal1 8142 29036 8142 29036 0 adapter.game.h\[4\]
rlabel metal1 23276 31926 23276 31926 0 adapter.game.h\[5\]
rlabel metal1 22908 32878 22908 32878 0 adapter.game.h\[6\]
rlabel metal1 18676 33830 18676 33830 0 adapter.game.h\[7\]
rlabel metal1 18722 34544 18722 34544 0 adapter.game.h\[8\]
rlabel metal2 17618 32572 17618 32572 0 adapter.game.h\[9\]
rlabel metal2 23322 16694 23322 16694 0 adapter.game.hit
rlabel metal1 4370 24650 4370 24650 0 adapter.game.hsync
rlabel metal1 24794 32402 24794 32402 0 adapter.game.inBallX
rlabel metal1 20470 20570 20470 20570 0 adapter.game.inBallY
rlabel metal1 16146 17034 16146 17034 0 adapter.game.inPaddle
rlabel metal1 19734 25670 19734 25670 0 adapter.game.offset\[0\]
rlabel metal1 15502 29070 15502 29070 0 adapter.game.offset\[1\]
rlabel metal2 14306 26180 14306 26180 0 adapter.game.offset\[2\]
rlabel metal1 12052 29818 12052 29818 0 adapter.game.offset\[3\]
rlabel metal1 8878 26962 8878 26962 0 adapter.game.offset\[4\]
rlabel metal1 15456 18598 15456 18598 0 adapter.game.paddle\[0\]
rlabel metal1 19412 15470 19412 15470 0 adapter.game.paddle\[1\]
rlabel metal1 18584 18326 18584 18326 0 adapter.game.paddle\[2\]
rlabel metal1 20424 14586 20424 14586 0 adapter.game.paddle\[3\]
rlabel metal1 20608 13974 20608 13974 0 adapter.game.paddle\[4\]
rlabel metal1 16698 13838 16698 13838 0 adapter.game.paddle\[5\]
rlabel metal1 13018 12716 13018 12716 0 adapter.game.paddle\[6\]
rlabel metal1 14812 12954 14812 12954 0 adapter.game.paddle\[7\]
rlabel metal1 14536 12886 14536 12886 0 adapter.game.paddle\[8\]
rlabel metal1 23322 34510 23322 34510 0 adapter.game.red
rlabel metal2 23828 16524 23828 16524 0 adapter.game.speaker
rlabel metal1 16008 19754 16008 19754 0 adapter.game.v\[0\]
rlabel metal1 15042 25262 15042 25262 0 adapter.game.v\[1\]
rlabel metal1 11776 24378 11776 24378 0 adapter.game.v\[2\]
rlabel metal1 12190 22984 12190 22984 0 adapter.game.v\[3\]
rlabel metal2 13018 21114 13018 21114 0 adapter.game.v\[4\]
rlabel metal2 13202 21658 13202 21658 0 adapter.game.v\[5\]
rlabel metal1 19550 19720 19550 19720 0 adapter.game.v\[6\]
rlabel metal2 13478 21216 13478 21216 0 adapter.game.v\[7\]
rlabel metal1 12098 18938 12098 18938 0 adapter.game.v\[8\]
rlabel metal1 14490 21522 14490 21522 0 adapter.game.v\[9\]
rlabel metal2 13754 24548 13754 24548 0 adapter.game.vsync
rlabel metal1 15686 18326 15686 18326 0 clknet_0_wb_clk_i
rlabel metal2 13846 17408 13846 17408 0 clknet_3_0__leaf_wb_clk_i
rlabel metal1 10764 23086 10764 23086 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 22034 16796 22034 16796 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 22034 20723 22034 20723 0 clknet_3_3__leaf_wb_clk_i
rlabel metal1 16790 32844 16790 32844 0 clknet_3_4__leaf_wb_clk_i
rlabel metal1 14812 35054 14812 35054 0 clknet_3_5__leaf_wb_clk_i
rlabel metal1 21528 26350 21528 26350 0 clknet_3_6__leaf_wb_clk_i
rlabel metal1 21666 33966 21666 33966 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 29026 1588 29026 1588 0 io_in[10]
rlabel metal2 30958 1554 30958 1554 0 io_in[11]
rlabel metal2 9062 1554 9062 1554 0 io_in[12]
rlabel metal3 1142 8228 1142 8228 0 io_in[8]
rlabel metal3 1188 3468 1188 3468 0 io_in[9]
rlabel metal2 26450 2166 26450 2166 0 io_oeb[0]
rlabel metal1 29624 36210 29624 36210 0 io_oeb[10]
rlabel metal2 34822 1860 34822 1860 0 io_oeb[11]
rlabel metal1 30360 37298 30360 37298 0 io_oeb[12]
rlabel metal2 35742 23817 35742 23817 0 io_oeb[13]
rlabel metal2 35742 31705 35742 31705 0 io_oeb[14]
rlabel metal2 35466 22389 35466 22389 0 io_oeb[15]
rlabel metal2 4094 12835 4094 12835 0 io_oeb[16]
rlabel metal1 19458 3366 19458 3366 0 io_oeb[17]
rlabel metal1 34776 34034 34776 34034 0 io_oeb[18]
rlabel metal3 1142 6868 1142 6868 0 io_oeb[19]
rlabel metal2 37122 3383 37122 3383 0 io_oeb[1]
rlabel metal3 1740 748 1740 748 0 io_oeb[20]
rlabel metal2 10994 2166 10994 2166 0 io_oeb[21]
rlabel metal3 37544 36788 37544 36788 0 io_oeb[22]
rlabel metal1 32798 36652 32798 36652 0 io_oeb[23]
rlabel metal2 3266 1231 3266 1231 0 io_oeb[24]
rlabel metal2 12282 1622 12282 1622 0 io_oeb[25]
rlabel metal2 37214 22287 37214 22287 0 io_oeb[26]
rlabel metal2 25162 1622 25162 1622 0 io_oeb[27]
rlabel via2 2806 12291 2806 12291 0 io_oeb[28]
rlabel metal2 18078 37954 18078 37954 0 io_oeb[29]
rlabel metal3 1142 29308 1142 29308 0 io_oeb[2]
rlabel metal1 4646 36652 4646 36652 0 io_oeb[30]
rlabel metal2 38686 38158 38686 38158 0 io_oeb[31]
rlabel metal2 22862 37349 22862 37349 0 io_oeb[32]
rlabel metal3 38786 34068 38786 34068 0 io_oeb[33]
rlabel metal2 37858 34935 37858 34935 0 io_oeb[34]
rlabel via2 4094 19805 4094 19805 0 io_oeb[35]
rlabel metal1 32936 37298 32936 37298 0 io_oeb[36]
rlabel metal2 37858 25279 37858 25279 0 io_oeb[37]
rlabel metal2 7130 37954 7130 37954 0 io_oeb[3]
rlabel metal2 37214 11067 37214 11067 0 io_oeb[4]
rlabel metal3 1740 33388 1740 33388 0 io_oeb[5]
rlabel metal1 4324 36210 4324 36210 0 io_oeb[6]
rlabel metal1 34224 37298 34224 37298 0 io_oeb[7]
rlabel metal2 37858 18955 37858 18955 0 io_oeb[8]
rlabel metal3 1280 17068 1280 17068 0 io_oeb[9]
rlabel metal3 1280 37468 1280 37468 0 io_out[0]
rlabel metal3 1786 1428 1786 1428 0 io_out[10]
rlabel metal2 21298 2166 21298 2166 0 io_out[11]
rlabel metal2 2806 17969 2806 17969 0 io_out[12]
rlabel metal2 24518 36866 24518 36866 0 io_out[13]
rlabel metal1 38594 37638 38594 37638 0 io_out[14]
rlabel metal1 4278 26418 4278 26418 0 io_out[15]
rlabel metal2 3910 2234 3910 2234 0 io_out[16]
rlabel metal1 15410 34714 15410 34714 0 io_out[17]
rlabel metal2 34546 9197 34546 9197 0 io_out[18]
rlabel metal2 34178 37551 34178 37551 0 io_out[19]
rlabel metal3 1832 2108 1832 2108 0 io_out[1]
rlabel metal2 2898 14943 2898 14943 0 io_out[20]
rlabel metal2 34178 1299 34178 1299 0 io_out[21]
rlabel metal2 37996 37604 37996 37604 0 io_out[22]
rlabel metal1 27646 36652 27646 36652 0 io_out[23]
rlabel metal2 37858 24395 37858 24395 0 io_out[24]
rlabel metal3 1878 29988 1878 29988 0 io_out[25]
rlabel metal2 39330 3288 39330 3288 0 io_out[26]
rlabel metal3 38786 17068 38786 17068 0 io_out[27]
rlabel metal2 23874 37920 23874 37920 0 io_out[28]
rlabel metal1 29854 36686 29854 36686 0 io_out[29]
rlabel metal2 37214 12631 37214 12631 0 io_out[2]
rlabel metal3 1878 2788 1878 2788 0 io_out[30]
rlabel metal2 25806 38260 25806 38260 0 io_out[31]
rlabel metal2 9706 37954 9706 37954 0 io_out[32]
rlabel metal2 16146 37716 16146 37716 0 io_out[33]
rlabel metal2 22080 36210 22080 36210 0 io_out[34]
rlabel metal2 38686 2098 38686 2098 0 io_out[35]
rlabel metal3 1142 8908 1142 8908 0 io_out[36]
rlabel metal2 35834 3417 35834 3417 0 io_out[37]
rlabel metal2 5842 3798 5842 3798 0 io_out[3]
rlabel metal2 2806 21947 2806 21947 0 io_out[4]
rlabel metal2 20654 37954 20654 37954 0 io_out[5]
rlabel metal3 38786 17748 38786 17748 0 io_out[6]
rlabel metal3 38234 7548 38234 7548 0 io_out[7]
rlabel metal2 2806 37179 2806 37179 0 io_out[8]
rlabel metal3 38786 33388 38786 33388 0 io_out[9]
rlabel metal1 2254 18632 2254 18632 0 net1
rlabel metal2 10626 27761 10626 27761 0 net10
rlabel metal1 22448 36686 22448 36686 0 net100
rlabel metal1 38134 33524 38134 33524 0 net101
rlabel metal2 38318 34816 38318 34816 0 net102
rlabel metal1 4324 28050 4324 28050 0 net103
rlabel metal1 32614 34442 32614 34442 0 net104
rlabel metal2 38318 25500 38318 25500 0 net105
rlabel metal2 2162 29580 2162 29580 0 net11
rlabel metal2 1886 14756 1886 14756 0 net12
rlabel metal1 27968 2618 27968 2618 0 net13
rlabel metal1 38088 7922 38088 7922 0 net14
rlabel via1 8234 4131 8234 4131 0 net15
rlabel metal2 12926 3264 12926 3264 0 net16
rlabel metal2 22034 3468 22034 3468 0 net17
rlabel metal2 36478 27676 36478 27676 0 net18
rlabel metal2 24334 3264 24334 3264 0 net19
rlabel metal1 29992 2482 29992 2482 0 net2
rlabel metal1 29072 35734 29072 35734 0 net20
rlabel metal1 27048 35258 27048 35258 0 net21
rlabel metal1 36478 15572 36478 15572 0 net22
rlabel metal2 8878 3264 8878 3264 0 net23
rlabel metal2 38318 30940 38318 30940 0 net24
rlabel metal2 37214 36380 37214 36380 0 net25
rlabel metal2 36938 3740 36938 3740 0 net26
rlabel metal1 34500 35258 34500 35258 0 net27
rlabel metal2 3082 20400 3082 20400 0 net28
rlabel metal2 3726 22848 3726 22848 0 net29
rlabel metal1 22540 2550 22540 2550 0 net3
rlabel metal2 5566 3740 5566 3740 0 net30
rlabel metal2 1886 5440 1886 5440 0 net31
rlabel metal2 1886 28288 1886 28288 0 net32
rlabel metal2 3910 32640 3910 32640 0 net33
rlabel metal2 18906 36720 18906 36720 0 net34
rlabel metal1 3634 20026 3634 20026 0 net35
rlabel metal1 6670 2618 6670 2618 0 net36
rlabel metal1 4324 2482 4324 2482 0 net37
rlabel metal1 24518 35666 24518 35666 0 net38
rlabel metal1 14720 36686 14720 36686 0 net39
rlabel metal1 10120 2414 10120 2414 0 net4
rlabel metal1 19504 3026 19504 3026 0 net40
rlabel metal1 31740 35666 31740 35666 0 net41
rlabel metal2 1610 31280 1610 31280 0 net42
rlabel metal1 38088 29138 38088 29138 0 net43
rlabel metal1 3726 36788 3726 36788 0 net44
rlabel metal1 3588 4046 3588 4046 0 net45
rlabel metal2 38318 12784 38318 12784 0 net46
rlabel metal2 5382 7004 5382 7004 0 net47
rlabel metal1 1656 21522 1656 21522 0 net48
rlabel metal1 19550 36754 19550 36754 0 net49
rlabel metal2 20470 17204 20470 17204 0 net5
rlabel metal2 36478 17884 36478 17884 0 net50
rlabel metal1 38088 8942 38088 8942 0 net51
rlabel metal1 1656 35666 1656 35666 0 net52
rlabel metal2 36478 33116 36478 33116 0 net53
rlabel metal1 4232 2958 4232 2958 0 net54
rlabel metal2 20746 3740 20746 3740 0 net55
rlabel metal1 1840 17850 1840 17850 0 net56
rlabel metal2 30038 3740 30038 3740 0 net57
rlabel metal1 37214 35598 37214 35598 0 net58
rlabel metal1 27186 36788 27186 36788 0 net59
rlabel via2 1886 2363 1886 2363 0 net6
rlabel metal2 38318 24412 38318 24412 0 net60
rlabel metal2 4094 30668 4094 30668 0 net61
rlabel metal1 38088 5202 38088 5202 0 net62
rlabel metal1 36478 16660 36478 16660 0 net63
rlabel metal1 24012 36754 24012 36754 0 net64
rlabel metal1 28980 36618 28980 36618 0 net65
rlabel metal1 2806 10574 2806 10574 0 net66
rlabel metal1 26910 37230 26910 37230 0 net67
rlabel metal2 9246 36992 9246 36992 0 net68
rlabel metal1 14628 36210 14628 36210 0 net69
rlabel metal2 38042 30481 38042 30481 0 net7
rlabel metal2 21022 36720 21022 36720 0 net70
rlabel metal2 36294 3298 36294 3298 0 net71
rlabel metal1 3450 9044 3450 9044 0 net72
rlabel metal1 37536 4046 37536 4046 0 net73
rlabel metal2 25898 4080 25898 4080 0 net74
rlabel metal1 38180 3026 38180 3026 0 net75
rlabel metal1 3220 29682 3220 29682 0 net76
rlabel metal2 6578 36992 6578 36992 0 net77
rlabel metal2 38318 11356 38318 11356 0 net78
rlabel metal2 1886 33728 1886 33728 0 net79
rlabel metal2 33902 28866 33902 28866 0 net8
rlabel metal1 3726 36210 3726 36210 0 net80
rlabel metal1 34960 34170 34960 34170 0 net81
rlabel metal2 38318 18972 38318 18972 0 net82
rlabel metal2 2162 16932 2162 16932 0 net83
rlabel metal1 29440 36142 29440 36142 0 net84
rlabel metal2 33994 3468 33994 3468 0 net85
rlabel metal1 30314 37094 30314 37094 0 net86
rlabel metal1 2806 7174 2806 7174 0 net87
rlabel metal1 3726 3570 3726 3570 0 net88
rlabel metal1 10212 3502 10212 3502 0 net89
rlabel metal2 33626 23936 33626 23936 0 net9
rlabel metal2 37674 33456 37674 33456 0 net90
rlabel metal2 32338 35972 32338 35972 0 net91
rlabel metal2 4186 3264 4186 3264 0 net92
rlabel metal2 11822 3196 11822 3196 0 net93
rlabel metal2 38318 22576 38318 22576 0 net94
rlabel metal2 24610 2992 24610 2992 0 net95
rlabel metal1 1748 11730 1748 11730 0 net96
rlabel metal2 19182 37026 19182 37026 0 net97
rlabel metal2 4186 36992 4186 36992 0 net98
rlabel metal1 36478 34170 36478 34170 0 net99
rlabel metal2 12604 39236 12604 39236 0 wb_clk_i
rlabel metal2 38318 38063 38318 38063 0 wb_rst_i
rlabel metal3 1786 28628 1786 28628 0 wbs_ack_o
rlabel metal2 2806 14977 2806 14977 0 wbs_dat_o[0]
rlabel metal3 38786 16388 38786 16388 0 wbs_dat_o[10]
rlabel metal2 690 1962 690 1962 0 wbs_dat_o[11]
rlabel metal2 37858 30719 37858 30719 0 wbs_dat_o[12]
rlabel metal1 36754 36244 36754 36244 0 wbs_dat_o[13]
rlabel metal1 36478 2516 36478 2516 0 wbs_dat_o[14]
rlabel metal2 34822 38277 34822 38277 0 wbs_dat_o[15]
rlabel metal3 1142 21148 1142 21148 0 wbs_dat_o[16]
rlabel metal3 1280 22508 1280 22508 0 wbs_dat_o[17]
rlabel metal2 24518 1299 24518 1299 0 wbs_dat_o[18]
rlabel metal2 46 2914 46 2914 0 wbs_dat_o[19]
rlabel metal2 28382 1860 28382 1860 0 wbs_dat_o[1]
rlabel metal3 1740 27948 1740 27948 0 wbs_dat_o[20]
rlabel metal2 2622 37551 2622 37551 0 wbs_dat_o[21]
rlabel metal2 17434 37716 17434 37716 0 wbs_dat_o[22]
rlabel metal3 1326 20468 1326 20468 0 wbs_dat_o[23]
rlabel metal2 7774 1860 7774 1860 0 wbs_dat_o[24]
rlabel metal2 2622 1792 2622 1792 0 wbs_dat_o[25]
rlabel metal2 25162 37716 25162 37716 0 wbs_dat_o[26]
rlabel metal2 16790 38022 16790 38022 0 wbs_dat_o[27]
rlabel metal2 20010 1860 20010 1860 0 wbs_dat_o[28]
rlabel metal1 31740 36210 31740 36210 0 wbs_dat_o[29]
rlabel metal2 37214 8075 37214 8075 0 wbs_dat_o[2]
rlabel metal3 1740 30668 1740 30668 0 wbs_dat_o[30]
rlabel metal2 37214 29155 37214 29155 0 wbs_dat_o[31]
rlabel metal2 8418 1503 8418 1503 0 wbs_dat_o[3]
rlabel metal2 13570 1860 13570 1860 0 wbs_dat_o[4]
rlabel metal2 22586 1860 22586 1860 0 wbs_dat_o[5]
rlabel metal3 38786 27268 38786 27268 0 wbs_dat_o[6]
rlabel metal2 23230 1826 23230 1826 0 wbs_dat_o[7]
rlabel metal1 27692 35734 27692 35734 0 wbs_dat_o[8]
rlabel metal1 27232 36210 27232 36210 0 wbs_dat_o[9]
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
