magic
tech sky130A
magscale 1 2
timestamp 1680612647
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37664
<< metal2 >>
rect -10 39200 102 39800
rect 634 39200 746 39800
rect 1278 39200 1390 39800
rect 1922 39200 2034 39800
rect 2566 39200 2678 39800
rect 3210 39200 3322 39800
rect 3854 39200 3966 39800
rect 4498 39200 4610 39800
rect 5142 39200 5254 39800
rect 5786 39200 5898 39800
rect 7074 39200 7186 39800
rect 7718 39200 7830 39800
rect 8362 39200 8474 39800
rect 9006 39200 9118 39800
rect 9650 39200 9762 39800
rect 10294 39200 10406 39800
rect 10938 39200 11050 39800
rect 11582 39200 11694 39800
rect 12226 39200 12338 39800
rect 12870 39200 12982 39800
rect 14158 39200 14270 39800
rect 14802 39200 14914 39800
rect 15446 39200 15558 39800
rect 16090 39200 16202 39800
rect 16734 39200 16846 39800
rect 17378 39200 17490 39800
rect 18022 39200 18134 39800
rect 18666 39200 18778 39800
rect 19310 39200 19422 39800
rect 19954 39200 20066 39800
rect 20598 39200 20710 39800
rect 21886 39200 21998 39800
rect 22530 39200 22642 39800
rect 23174 39200 23286 39800
rect 23818 39200 23930 39800
rect 24462 39200 24574 39800
rect 25106 39200 25218 39800
rect 25750 39200 25862 39800
rect 26394 39200 26506 39800
rect 27038 39200 27150 39800
rect 27682 39200 27794 39800
rect 28970 39200 29082 39800
rect 29614 39200 29726 39800
rect 30258 39200 30370 39800
rect 30902 39200 31014 39800
rect 31546 39200 31658 39800
rect 32190 39200 32302 39800
rect 32834 39200 32946 39800
rect 33478 39200 33590 39800
rect 34122 39200 34234 39800
rect 34766 39200 34878 39800
rect 35410 39200 35522 39800
rect 36698 39200 36810 39800
rect 37342 39200 37454 39800
rect 37986 39200 38098 39800
rect 38630 39200 38742 39800
rect 39274 39200 39386 39800
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5142 200 5254 800
rect 5786 200 5898 800
rect 6430 200 6542 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10294 200 10406 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12226 200 12338 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 15446 200 15558 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 18666 200 18778 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 20598 200 20710 800
rect 21242 200 21354 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25106 200 25218 800
rect 25750 200 25862 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 30258 200 30370 800
rect 30902 200 31014 800
rect 31546 200 31658 800
rect 32190 200 32302 800
rect 32834 200 32946 800
rect 33478 200 33590 800
rect 34122 200 34234 800
rect 34766 200 34878 800
rect 35410 200 35522 800
rect 36054 200 36166 800
rect 37342 200 37454 800
rect 37986 200 38098 800
rect 38630 200 38742 800
rect 39274 200 39386 800
<< obsm2 >>
rect 158 39144 578 39250
rect 802 39144 1222 39250
rect 1446 39144 1866 39250
rect 2090 39144 2510 39250
rect 2734 39144 3154 39250
rect 3378 39144 3798 39250
rect 4022 39144 4442 39250
rect 4666 39144 5086 39250
rect 5310 39144 5730 39250
rect 5954 39144 7018 39250
rect 7242 39144 7662 39250
rect 7886 39144 8306 39250
rect 8530 39144 8950 39250
rect 9174 39144 9594 39250
rect 9818 39144 10238 39250
rect 10462 39144 10882 39250
rect 11106 39144 11526 39250
rect 11750 39144 12170 39250
rect 12394 39144 12814 39250
rect 13038 39144 14102 39250
rect 14326 39144 14746 39250
rect 14970 39144 15390 39250
rect 15614 39144 16034 39250
rect 16258 39144 16678 39250
rect 16902 39144 17322 39250
rect 17546 39144 17966 39250
rect 18190 39144 18610 39250
rect 18834 39144 19254 39250
rect 19478 39144 19898 39250
rect 20122 39144 20542 39250
rect 20766 39144 21830 39250
rect 22054 39144 22474 39250
rect 22698 39144 23118 39250
rect 23342 39144 23762 39250
rect 23986 39144 24406 39250
rect 24630 39144 25050 39250
rect 25274 39144 25694 39250
rect 25918 39144 26338 39250
rect 26562 39144 26982 39250
rect 27206 39144 27626 39250
rect 27850 39144 28914 39250
rect 29138 39144 29558 39250
rect 29782 39144 30202 39250
rect 30426 39144 30846 39250
rect 31070 39144 31490 39250
rect 31714 39144 32134 39250
rect 32358 39144 32778 39250
rect 33002 39144 33422 39250
rect 33646 39144 34066 39250
rect 34290 39144 34710 39250
rect 34934 39144 35354 39250
rect 35578 39144 36642 39250
rect 36866 39144 37286 39250
rect 37510 39144 37930 39250
rect 38154 39144 38574 39250
rect 38798 39144 39218 39250
rect 20 856 39356 39144
rect 158 144 578 856
rect 802 144 1222 856
rect 1446 144 1866 856
rect 2090 144 2510 856
rect 2734 144 3154 856
rect 3378 144 3798 856
rect 4022 144 4442 856
rect 4666 144 5086 856
rect 5310 144 5730 856
rect 5954 144 6374 856
rect 6598 144 7662 856
rect 7886 144 8306 856
rect 8530 144 8950 856
rect 9174 144 9594 856
rect 9818 144 10238 856
rect 10462 144 10882 856
rect 11106 144 11526 856
rect 11750 144 12170 856
rect 12394 144 12814 856
rect 13038 144 13458 856
rect 13682 144 14102 856
rect 14326 144 15390 856
rect 15614 144 16034 856
rect 16258 144 16678 856
rect 16902 144 17322 856
rect 17546 144 17966 856
rect 18190 144 18610 856
rect 18834 144 19254 856
rect 19478 144 19898 856
rect 20122 144 20542 856
rect 20766 144 21186 856
rect 21410 144 22474 856
rect 22698 144 23118 856
rect 23342 144 23762 856
rect 23986 144 24406 856
rect 24630 144 25050 856
rect 25274 144 25694 856
rect 25918 144 26338 856
rect 26562 144 26982 856
rect 27206 144 27626 856
rect 27850 144 28270 856
rect 28494 144 28914 856
rect 29138 144 30202 856
rect 30426 144 30846 856
rect 31070 144 31490 856
rect 31714 144 32134 856
rect 32358 144 32778 856
rect 33002 144 33422 856
rect 33646 144 34066 856
rect 34290 144 34710 856
rect 34934 144 35354 856
rect 35578 144 35998 856
rect 36222 144 37286 856
rect 37510 144 37930 856
rect 38154 144 38574 856
rect 38798 144 39218 856
rect 20 31 39356 144
<< metal3 >>
rect 200 39388 800 39628
rect 39200 39388 39800 39628
rect 39200 38708 39800 38948
rect 200 38028 800 38268
rect 39200 38028 39800 38268
rect 200 37348 800 37588
rect 39200 37348 39800 37588
rect 200 36668 800 36908
rect 39200 36668 39800 36908
rect 200 35988 800 36228
rect 200 35308 800 35548
rect 39200 35308 39800 35548
rect 200 34628 800 34868
rect 39200 34628 39800 34868
rect 200 33948 800 34188
rect 39200 33948 39800 34188
rect 200 33268 800 33508
rect 39200 33268 39800 33508
rect 200 32588 800 32828
rect 39200 32588 39800 32828
rect 200 31908 800 32148
rect 39200 31908 39800 32148
rect 39200 31228 39800 31468
rect 200 30548 800 30788
rect 39200 30548 39800 30788
rect 200 29868 800 30108
rect 39200 29868 39800 30108
rect 200 29188 800 29428
rect 39200 29188 39800 29428
rect 200 28508 800 28748
rect 39200 28508 39800 28748
rect 200 27828 800 28068
rect 200 27148 800 27388
rect 39200 27148 39800 27388
rect 200 26468 800 26708
rect 39200 26468 39800 26708
rect 200 25788 800 26028
rect 39200 25788 39800 26028
rect 200 25108 800 25348
rect 39200 25108 39800 25348
rect 200 24428 800 24668
rect 39200 24428 39800 24668
rect 200 23748 800 23988
rect 39200 23748 39800 23988
rect 39200 23068 39800 23308
rect 200 22388 800 22628
rect 39200 22388 39800 22628
rect 200 21708 800 21948
rect 39200 21708 39800 21948
rect 200 21028 800 21268
rect 39200 21028 39800 21268
rect 200 20348 800 20588
rect 200 19668 800 19908
rect 39200 19668 39800 19908
rect 200 18988 800 19228
rect 39200 18988 39800 19228
rect 200 18308 800 18548
rect 39200 18308 39800 18548
rect 200 17628 800 17868
rect 39200 17628 39800 17868
rect 200 16948 800 17188
rect 39200 16948 39800 17188
rect 200 16268 800 16508
rect 39200 16268 39800 16508
rect 39200 15588 39800 15828
rect 200 14908 800 15148
rect 39200 14908 39800 15148
rect 200 14228 800 14468
rect 39200 14228 39800 14468
rect 200 13548 800 13788
rect 39200 13548 39800 13788
rect 200 12868 800 13108
rect 39200 12868 39800 13108
rect 200 12188 800 12428
rect 200 11508 800 11748
rect 39200 11508 39800 11748
rect 200 10828 800 11068
rect 39200 10828 39800 11068
rect 200 10148 800 10388
rect 39200 10148 39800 10388
rect 200 9468 800 9708
rect 39200 9468 39800 9708
rect 200 8788 800 9028
rect 39200 8788 39800 9028
rect 200 8108 800 8348
rect 39200 8108 39800 8348
rect 39200 7428 39800 7668
rect 200 6748 800 6988
rect 39200 6748 39800 6988
rect 200 6068 800 6308
rect 39200 6068 39800 6308
rect 200 5388 800 5628
rect 39200 5388 39800 5628
rect 200 4708 800 4948
rect 200 4028 800 4268
rect 39200 4028 39800 4268
rect 200 3348 800 3588
rect 39200 3348 39800 3588
rect 200 2668 800 2908
rect 39200 2668 39800 2908
rect 200 1988 800 2228
rect 39200 1988 39800 2228
rect 200 1308 800 1548
rect 39200 1308 39800 1548
rect 200 628 800 868
rect 39200 628 39800 868
rect 39200 -52 39800 188
<< obsm3 >>
rect 800 38628 39120 38861
rect 800 38348 39200 38628
rect 880 37948 39120 38348
rect 800 37668 39200 37948
rect 880 37268 39120 37668
rect 800 36988 39200 37268
rect 880 36588 39120 36988
rect 800 36308 39200 36588
rect 880 35908 39200 36308
rect 800 35628 39200 35908
rect 880 35228 39120 35628
rect 800 34948 39200 35228
rect 880 34548 39120 34948
rect 800 34268 39200 34548
rect 880 33868 39120 34268
rect 800 33588 39200 33868
rect 880 33188 39120 33588
rect 800 32908 39200 33188
rect 880 32508 39120 32908
rect 800 32228 39200 32508
rect 880 31828 39120 32228
rect 800 31548 39200 31828
rect 800 31148 39120 31548
rect 800 30868 39200 31148
rect 880 30468 39120 30868
rect 800 30188 39200 30468
rect 880 29788 39120 30188
rect 800 29508 39200 29788
rect 880 29108 39120 29508
rect 800 28828 39200 29108
rect 880 28428 39120 28828
rect 800 28148 39200 28428
rect 880 27748 39200 28148
rect 800 27468 39200 27748
rect 880 27068 39120 27468
rect 800 26788 39200 27068
rect 880 26388 39120 26788
rect 800 26108 39200 26388
rect 880 25708 39120 26108
rect 800 25428 39200 25708
rect 880 25028 39120 25428
rect 800 24748 39200 25028
rect 880 24348 39120 24748
rect 800 24068 39200 24348
rect 880 23668 39120 24068
rect 800 23388 39200 23668
rect 800 22988 39120 23388
rect 800 22708 39200 22988
rect 880 22308 39120 22708
rect 800 22028 39200 22308
rect 880 21628 39120 22028
rect 800 21348 39200 21628
rect 880 20948 39120 21348
rect 800 20668 39200 20948
rect 880 20268 39200 20668
rect 800 19988 39200 20268
rect 880 19588 39120 19988
rect 800 19308 39200 19588
rect 880 18908 39120 19308
rect 800 18628 39200 18908
rect 880 18228 39120 18628
rect 800 17948 39200 18228
rect 880 17548 39120 17948
rect 800 17268 39200 17548
rect 880 16868 39120 17268
rect 800 16588 39200 16868
rect 880 16188 39120 16588
rect 800 15908 39200 16188
rect 800 15508 39120 15908
rect 800 15228 39200 15508
rect 880 14828 39120 15228
rect 800 14548 39200 14828
rect 880 14148 39120 14548
rect 800 13868 39200 14148
rect 880 13468 39120 13868
rect 800 13188 39200 13468
rect 880 12788 39120 13188
rect 800 12508 39200 12788
rect 880 12108 39200 12508
rect 800 11828 39200 12108
rect 880 11428 39120 11828
rect 800 11148 39200 11428
rect 880 10748 39120 11148
rect 800 10468 39200 10748
rect 880 10068 39120 10468
rect 800 9788 39200 10068
rect 880 9388 39120 9788
rect 800 9108 39200 9388
rect 880 8708 39120 9108
rect 800 8428 39200 8708
rect 880 8028 39120 8428
rect 800 7748 39200 8028
rect 800 7348 39120 7748
rect 800 7068 39200 7348
rect 880 6668 39120 7068
rect 800 6388 39200 6668
rect 880 5988 39120 6388
rect 800 5708 39200 5988
rect 880 5308 39120 5708
rect 800 5028 39200 5308
rect 880 4628 39200 5028
rect 800 4348 39200 4628
rect 880 3948 39120 4348
rect 800 3668 39200 3948
rect 880 3268 39120 3668
rect 800 2988 39200 3268
rect 880 2588 39120 2988
rect 800 2308 39200 2588
rect 880 1908 39120 2308
rect 800 1628 39200 1908
rect 880 1228 39120 1628
rect 800 948 39200 1228
rect 880 548 39120 948
rect 800 268 39200 548
rect 800 35 39120 268
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 17355 2347 17421 20909
<< labels >>
rlabel metal2 s -10 39200 102 39800 6 active
port 1 nsew signal input
rlabel metal3 s 39200 11508 39800 11748 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 28970 200 29082 800 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 30902 200 31014 800 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 9006 200 9118 800 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 39200 6068 39800 6308 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 39200 4028 39800 4268 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 14158 200 14270 800 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 200 5388 800 5628 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 39200 19668 39800 19908 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 39200 14908 39800 15148 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 32190 200 32302 800 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 12226 39200 12338 39800 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 39200 628 39800 868 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 39200 29188 39800 29428 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 5142 39200 5254 39800 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 33478 39200 33590 39800 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 200 27148 800 27388 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 36698 39200 36810 39800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 18666 39200 18778 39800 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 30258 200 30370 800 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 200 4708 800 4948 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 25750 200 25862 800 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 7718 39200 7830 39800 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 1278 39200 1390 39800 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 10294 39200 10406 39800 6 io_in[31]
port 26 nsew signal input
rlabel metal3 s 200 16268 800 16508 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 39200 1308 39800 1548 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 20598 200 20710 800 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 39200 13548 39800 13788 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 200 35988 800 36228 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 39200 26468 39800 26708 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 33478 200 33590 800 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 200 32588 800 32828 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 12870 200 12982 800 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 17378 200 17490 800 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 32834 200 32946 800 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 200 8108 800 8348 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 200 3348 800 3588 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 26394 200 26506 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal2 s 28970 39200 29082 39800 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal2 s 34766 200 34878 800 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal2 s 30258 39200 30370 39800 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal3 s 39200 23748 39800 23988 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 39200 31908 39800 32148 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal3 s 39200 23068 39800 23308 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal3 s 200 12868 800 13108 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal2 s 19310 200 19422 800 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 35410 39200 35522 39800 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal3 s 200 6748 800 6988 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal3 s 39200 1988 39800 2228 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 200 628 800 868 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 10938 200 11050 800 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal3 s 39200 36668 39800 36908 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 32190 39200 32302 39800 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 3210 200 3322 800 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal2 s 12226 200 12338 800 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 39200 22388 39800 22628 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal2 s 25106 200 25218 800 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal3 s 200 12188 800 12428 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal2 s 18022 39200 18134 39800 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal3 s 200 29188 800 29428 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal2 s 3210 39200 3322 39800 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 38630 39200 38742 39800 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal2 s 22530 39200 22642 39800 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal3 s 39200 33948 39800 34188 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal3 s 39200 34628 39800 34868 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 200 19668 800 19908 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal2 s 32834 39200 32946 39800 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 39200 25108 39800 25348 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal2 s 7074 39200 7186 39800 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 39200 10828 39800 11068 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 200 33268 800 33508 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal2 s 3854 39200 3966 39800 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 39200 37348 39800 37588 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal3 s 39200 18988 39800 19228 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal3 s 200 16948 800 17188 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal3 s 200 37348 800 37588 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 200 1308 800 1548 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal2 s 21242 200 21354 800 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 200 17628 800 17868 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal2 s 24462 39200 24574 39800 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal2 s 39274 39200 39386 39800 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 200 26468 800 26708 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal2 s 3854 200 3966 800 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 14802 39200 14914 39800 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal3 s 39200 8788 39800 9028 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal2 s 34122 39200 34234 39800 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal3 s 200 1988 800 2228 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal3 s 200 14228 800 14468 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal2 s 34122 200 34234 800 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal2 s 37986 39200 38098 39800 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal2 s 26394 39200 26506 39800 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 39200 24428 39800 24668 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal3 s 200 29868 800 30108 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal2 s 39274 200 39386 800 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal3 s 39200 16948 39800 17188 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 23818 39200 23930 39800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal2 s 29614 39200 29726 39800 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal3 s 39200 12868 39800 13108 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 200 2668 800 2908 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal2 s 25750 39200 25862 39800 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal2 s 9650 39200 9762 39800 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal2 s 16090 39200 16202 39800 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal2 s 21886 39200 21998 39800 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal2 s 38630 200 38742 800 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal3 s 200 8788 800 9028 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal3 s 39200 2668 39800 2908 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal2 s 5786 200 5898 800 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal3 s 200 21708 800 21948 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 20598 39200 20710 39800 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal3 s 39200 17628 39800 17868 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 39200 7428 39800 7668 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal3 s 200 38028 800 38268 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 39200 33268 39800 33508 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 116 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 117 nsew ground bidirectional
rlabel metal2 s 12870 39200 12982 39800 6 wb_clk_i
port 118 nsew signal input
rlabel metal3 s 39200 38708 39800 38948 6 wb_rst_i
port 119 nsew signal input
rlabel metal3 s 200 28508 800 28748 6 wbs_ack_o
port 120 nsew signal bidirectional
rlabel metal3 s 39200 25788 39800 26028 6 wbs_adr_i[0]
port 121 nsew signal input
rlabel metal3 s 39200 32588 39800 32828 6 wbs_adr_i[10]
port 122 nsew signal input
rlabel metal3 s 200 23748 800 23988 6 wbs_adr_i[11]
port 123 nsew signal input
rlabel metal2 s 1922 200 2034 800 6 wbs_adr_i[12]
port 124 nsew signal input
rlabel metal2 s 15446 200 15558 800 6 wbs_adr_i[13]
port 125 nsew signal input
rlabel metal3 s 39200 9468 39800 9708 6 wbs_adr_i[14]
port 126 nsew signal input
rlabel metal2 s 19954 39200 20066 39800 6 wbs_adr_i[15]
port 127 nsew signal input
rlabel metal2 s 18022 200 18134 800 6 wbs_adr_i[16]
port 128 nsew signal input
rlabel metal3 s 39200 6748 39800 6988 6 wbs_adr_i[17]
port 129 nsew signal input
rlabel metal2 s 37986 200 38098 800 6 wbs_adr_i[18]
port 130 nsew signal input
rlabel metal3 s 200 35308 800 35548 6 wbs_adr_i[19]
port 131 nsew signal input
rlabel metal3 s 200 25788 800 26028 6 wbs_adr_i[1]
port 132 nsew signal input
rlabel metal3 s 39200 21708 39800 21948 6 wbs_adr_i[20]
port 133 nsew signal input
rlabel metal3 s 200 31908 800 32148 6 wbs_adr_i[21]
port 134 nsew signal input
rlabel metal3 s 200 13548 800 13788 6 wbs_adr_i[22]
port 135 nsew signal input
rlabel metal2 s 36054 200 36166 800 6 wbs_adr_i[23]
port 136 nsew signal input
rlabel metal2 s 11582 39200 11694 39800 6 wbs_adr_i[24]
port 137 nsew signal input
rlabel metal2 s 16090 200 16202 800 6 wbs_adr_i[25]
port 138 nsew signal input
rlabel metal3 s 200 18988 800 19228 6 wbs_adr_i[26]
port 139 nsew signal input
rlabel metal3 s 200 25108 800 25348 6 wbs_adr_i[27]
port 140 nsew signal input
rlabel metal3 s 200 11508 800 11748 6 wbs_adr_i[28]
port 141 nsew signal input
rlabel metal2 s 10938 39200 11050 39800 6 wbs_adr_i[29]
port 142 nsew signal input
rlabel metal2 s 11582 200 11694 800 6 wbs_adr_i[2]
port 143 nsew signal input
rlabel metal2 s 4498 39200 4610 39800 6 wbs_adr_i[30]
port 144 nsew signal input
rlabel metal3 s 39200 3348 39800 3588 6 wbs_adr_i[31]
port 145 nsew signal input
rlabel metal2 s 23818 200 23930 800 6 wbs_adr_i[3]
port 146 nsew signal input
rlabel metal3 s 39200 31228 39800 31468 6 wbs_adr_i[4]
port 147 nsew signal input
rlabel metal3 s 200 4028 800 4268 6 wbs_adr_i[5]
port 148 nsew signal input
rlabel metal2 s 9650 200 9762 800 6 wbs_adr_i[6]
port 149 nsew signal input
rlabel metal2 s 8362 39200 8474 39800 6 wbs_adr_i[7]
port 150 nsew signal input
rlabel metal2 s 31546 200 31658 800 6 wbs_adr_i[8]
port 151 nsew signal input
rlabel metal3 s 200 24428 800 24668 6 wbs_adr_i[9]
port 152 nsew signal input
rlabel metal2 s 31546 39200 31658 39800 6 wbs_cyc_i
port 153 nsew signal input
rlabel metal2 s 634 39200 746 39800 6 wbs_dat_i[0]
port 154 nsew signal input
rlabel metal2 s 9006 39200 9118 39800 6 wbs_dat_i[10]
port 155 nsew signal input
rlabel metal2 s 15446 39200 15558 39800 6 wbs_dat_i[11]
port 156 nsew signal input
rlabel metal2 s 14158 39200 14270 39800 6 wbs_dat_i[12]
port 157 nsew signal input
rlabel metal2 s 1278 200 1390 800 6 wbs_dat_i[13]
port 158 nsew signal input
rlabel metal2 s 6430 200 6542 800 6 wbs_dat_i[14]
port 159 nsew signal input
rlabel metal3 s 200 10828 800 11068 6 wbs_dat_i[15]
port 160 nsew signal input
rlabel metal2 s 18666 200 18778 800 6 wbs_dat_i[16]
port 161 nsew signal input
rlabel metal3 s 39200 38028 39800 38268 6 wbs_dat_i[17]
port 162 nsew signal input
rlabel metal2 s 1922 39200 2034 39800 6 wbs_dat_i[18]
port 163 nsew signal input
rlabel metal2 s 19310 39200 19422 39800 6 wbs_dat_i[19]
port 164 nsew signal input
rlabel metal2 s 4498 200 4610 800 6 wbs_dat_i[1]
port 165 nsew signal input
rlabel metal3 s 39200 14228 39800 14468 6 wbs_dat_i[20]
port 166 nsew signal input
rlabel metal3 s 39200 29868 39800 30108 6 wbs_dat_i[21]
port 167 nsew signal input
rlabel metal3 s 200 18308 800 18548 6 wbs_dat_i[22]
port 168 nsew signal input
rlabel metal3 s 39200 21028 39800 21268 6 wbs_dat_i[23]
port 169 nsew signal input
rlabel metal3 s 200 34628 800 34868 6 wbs_dat_i[24]
port 170 nsew signal input
rlabel metal3 s 200 6068 800 6308 6 wbs_dat_i[25]
port 171 nsew signal input
rlabel metal3 s 39200 35308 39800 35548 6 wbs_dat_i[26]
port 172 nsew signal input
rlabel metal2 s 23174 39200 23286 39800 6 wbs_dat_i[27]
port 173 nsew signal input
rlabel metal2 s 10294 200 10406 800 6 wbs_dat_i[28]
port 174 nsew signal input
rlabel metal3 s 39200 15588 39800 15828 6 wbs_dat_i[29]
port 175 nsew signal input
rlabel metal2 s 27682 200 27794 800 6 wbs_dat_i[2]
port 176 nsew signal input
rlabel metal3 s 39200 5388 39800 5628 6 wbs_dat_i[30]
port 177 nsew signal input
rlabel metal3 s 200 36668 800 36908 6 wbs_dat_i[31]
port 178 nsew signal input
rlabel metal2 s 35410 200 35522 800 6 wbs_dat_i[3]
port 179 nsew signal input
rlabel metal2 s 5142 200 5254 800 6 wbs_dat_i[4]
port 180 nsew signal input
rlabel metal2 s 16734 200 16846 800 6 wbs_dat_i[5]
port 181 nsew signal input
rlabel metal3 s 39200 10148 39800 10388 6 wbs_dat_i[6]
port 182 nsew signal input
rlabel metal3 s 39200 39388 39800 39628 6 wbs_dat_i[7]
port 183 nsew signal input
rlabel metal3 s 200 10148 800 10388 6 wbs_dat_i[8]
port 184 nsew signal input
rlabel metal2 s 37342 200 37454 800 6 wbs_dat_i[9]
port 185 nsew signal input
rlabel metal3 s 200 14908 800 15148 6 wbs_dat_o[0]
port 186 nsew signal bidirectional
rlabel metal3 s 39200 16268 39800 16508 6 wbs_dat_o[10]
port 187 nsew signal bidirectional
rlabel metal2 s 634 200 746 800 6 wbs_dat_o[11]
port 188 nsew signal bidirectional
rlabel metal3 s 39200 30548 39800 30788 6 wbs_dat_o[12]
port 189 nsew signal bidirectional
rlabel metal2 s 37342 39200 37454 39800 6 wbs_dat_o[13]
port 190 nsew signal bidirectional
rlabel metal3 s 39200 -52 39800 188 6 wbs_dat_o[14]
port 191 nsew signal bidirectional
rlabel metal2 s 34766 39200 34878 39800 6 wbs_dat_o[15]
port 192 nsew signal bidirectional
rlabel metal3 s 200 21028 800 21268 6 wbs_dat_o[16]
port 193 nsew signal bidirectional
rlabel metal3 s 200 22388 800 22628 6 wbs_dat_o[17]
port 194 nsew signal bidirectional
rlabel metal2 s 24462 200 24574 800 6 wbs_dat_o[18]
port 195 nsew signal bidirectional
rlabel metal2 s -10 200 102 800 6 wbs_dat_o[19]
port 196 nsew signal bidirectional
rlabel metal2 s 28326 200 28438 800 6 wbs_dat_o[1]
port 197 nsew signal bidirectional
rlabel metal3 s 200 27828 800 28068 6 wbs_dat_o[20]
port 198 nsew signal bidirectional
rlabel metal2 s 2566 39200 2678 39800 6 wbs_dat_o[21]
port 199 nsew signal bidirectional
rlabel metal2 s 17378 39200 17490 39800 6 wbs_dat_o[22]
port 200 nsew signal bidirectional
rlabel metal3 s 200 20348 800 20588 6 wbs_dat_o[23]
port 201 nsew signal bidirectional
rlabel metal2 s 7718 200 7830 800 6 wbs_dat_o[24]
port 202 nsew signal bidirectional
rlabel metal2 s 2566 200 2678 800 6 wbs_dat_o[25]
port 203 nsew signal bidirectional
rlabel metal2 s 25106 39200 25218 39800 6 wbs_dat_o[26]
port 204 nsew signal bidirectional
rlabel metal2 s 16734 39200 16846 39800 6 wbs_dat_o[27]
port 205 nsew signal bidirectional
rlabel metal2 s 19954 200 20066 800 6 wbs_dat_o[28]
port 206 nsew signal bidirectional
rlabel metal2 s 30902 39200 31014 39800 6 wbs_dat_o[29]
port 207 nsew signal bidirectional
rlabel metal3 s 39200 8108 39800 8348 6 wbs_dat_o[2]
port 208 nsew signal bidirectional
rlabel metal3 s 200 30548 800 30788 6 wbs_dat_o[30]
port 209 nsew signal bidirectional
rlabel metal3 s 39200 28508 39800 28748 6 wbs_dat_o[31]
port 210 nsew signal bidirectional
rlabel metal2 s 8362 200 8474 800 6 wbs_dat_o[3]
port 211 nsew signal bidirectional
rlabel metal2 s 13514 200 13626 800 6 wbs_dat_o[4]
port 212 nsew signal bidirectional
rlabel metal2 s 22530 200 22642 800 6 wbs_dat_o[5]
port 213 nsew signal bidirectional
rlabel metal3 s 39200 27148 39800 27388 6 wbs_dat_o[6]
port 214 nsew signal bidirectional
rlabel metal2 s 23174 200 23286 800 6 wbs_dat_o[7]
port 215 nsew signal bidirectional
rlabel metal2 s 27682 39200 27794 39800 6 wbs_dat_o[8]
port 216 nsew signal bidirectional
rlabel metal2 s 27038 39200 27150 39800 6 wbs_dat_o[9]
port 217 nsew signal bidirectional
rlabel metal3 s 200 39388 800 39628 6 wbs_sel_i[0]
port 218 nsew signal input
rlabel metal2 s 5786 39200 5898 39800 6 wbs_sel_i[1]
port 219 nsew signal input
rlabel metal2 s 27038 200 27150 800 6 wbs_sel_i[2]
port 220 nsew signal input
rlabel metal3 s 200 9468 800 9708 6 wbs_sel_i[3]
port 221 nsew signal input
rlabel metal3 s 200 33948 800 34188 6 wbs_stb_i
port 222 nsew signal input
rlabel metal3 s 39200 18308 39800 18548 6 wbs_we_i
port 223 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2548086
string GDS_FILE /openlane/designs/wrapped_solo_squash/runs/RUN_2023.04.04_12.47.15/results/signoff/wrapped_solo_squash.magic.gds
string GDS_START 427740
<< end >>

